
.SUBCKT PIPO_and_Combinational clk rst xin0 xin1 xin2 xin3 yin0 yin1 yin2 yin3 vddio r_out vdd vss


c1 vdd vss 1.05148e-15
c2 clk vss 169.772e-18
c3 rst vss 208.837e-18
c4 r_out vss 36.4081e-18
c5 vddio vss 49.3446e-18
c6 xin0 vss 47.6761e-18
c7 xin1 vss 53.9727e-18
c8 xin2 vss 57.9603e-18
c9 xin3 vss 60.8749e-18
c10 yin0 vss 43.5999e-18
c11 yin1 vss 49.5315e-18
c12 yin2 vss 51.5228e-18
c13 yin3 vss 60.2306e-18
c14 clk4 vss 27.1014e-18
c15 clk4b vss 95.3554e-18
c16 clkb vss 216.414e-18
c17 clk2 vss 25.8153e-18
c18 x0 vss 40.1396e-18
c19 x1 vss 40.2644e-18
c20 x2 vss 44.6484e-18
c21 x3 vss 47.1718e-18
c22 y0 vss 53.7371e-18
c23 y1 vss 53.4488e-18
c24 y2 vss 55.5271e-18
c25 y3 vss 55.321e-18
c26 net12 vss 92.2494e-18
c27 c1 vss 51.9719e-18
c28 c0 vss 51.689e-18
c29 r2 vss 74.4362e-18
c30 r1 vss 68.8447e-18
c31 a0 vss 104.934e-18
c32 a1 vss 55.9119e-18
c33 s0 vss 50.178e-18
c34 s1 vss 56.6335e-18
c35 r0 vss 141.399e-18
c36 a2 vss 103.688e-18
c37 a3 vss 55.4149e-18
c38 serial_out vss 105.736e-18
c39 i12__net3 vss 59.6419e-18
c40 i6__net3 vss 129.969e-18
c41 net5 vss 112.682e-18
c42 r_in vss 108.714e-18
c43 i12__net1 vss 62.8924e-18
c44 i12__net2 vss 58.5464e-18
c45 i11__net1 vss 108.186e-18
c46 i6__net2 vss 110.307e-18
c47 i6__abar vss 69.1677e-18
c48 i6__net4 vss 95.9298e-18
c49 i6__bbar vss 65.3991e-18
c50 i6__net1 vss 117.199e-18
c51 i5__net3 vss 135.29e-18
c52 i5__net2 vss 107.96e-18
c53 i5__abar vss 68.4173e-18
c54 i5__net4 vss 95.2949e-18
c55 i5__bbar vss 67.3721e-18
c56 i5__net1 vss 108.097e-18
c57 i4__net3 vss 121.614e-18
c58 i4__net2 vss 112.075e-18
c59 i4__abar vss 67.6781e-18
c60 i4__net4 vss 95.3001e-18
c61 i4__bbar vss 66.0874e-18
c62 i4__net1 vss 111.112e-18
c63 i3__net3 vss 121.249e-18
c64 i3__net2 vss 110.488e-18
c65 i3__abar vss 68.2929e-18
c66 i3__net4 vss 94.8226e-18
c67 i3__bbar vss 67.0316e-18
c68 i3__net1 vss 108.836e-18
c69 i14__i5__net3 vss 76.6851e-18
c70 i14__i5__net4 vss 98.5202e-18
c71 i14__i5__net5 vss 54.5552e-18
c72 i14__i5__net2 vss 79.2728e-18
c73 i14__i5__net1 vss 105.925e-18
c74 i14__i5__rstb vss 27.385e-18
c75 i14__i4__net3 vss 83.0685e-18
c76 i14__i4__net4 vss 98.4859e-18
c77 i14__i4__net5 vss 54.1774e-18
c78 i14__i4__net2 vss 77.8714e-18
c79 i14__i4__net1 vss 108.483e-18
c80 i14__net15 vss 59.0727e-18
c81 i14__i4__rstb vss 27.5166e-18
c82 i14__i3__net3 vss 82.9195e-18
c83 i14__i3__net4 vss 98.5002e-18
c84 i14__i3__net5 vss 54.4651e-18
c85 i14__i3__net2 vss 77.5308e-18
c86 i14__i3__net1 vss 108.614e-18
c87 i14__net9 vss 58.8515e-18
c88 i14__i3__rstb vss 27.5366e-18
c89 i14__i7__net2 vss 105.666e-18
c90 i14__net14 vss 131.807e-18
c91 i14__i2__net1 vss 33.145e-18
c92 i14__i1__net1 vss 33.0593e-18
c93 i14__net8 vss 129.993e-18
c94 i14__net2 vss 181.644e-18
c95 i14__i0__net1 vss 32.3656e-18
c96 i14__shift vss 33.3836e-18
c97 i14__i7__net1 vss 24.9123e-18
c98 i8__net1 vss 88.8747e-18
c99 i8__carry_bar vss 44.4402e-18
c100 i8__net49 vss 121.717e-18
c101 i8__net51 vss 58.2722e-18
c102 i8__net50 vss 97.7847e-18
c103 i8__net52 vss 103.673e-18
c104 i9__net1 vss 84.7298e-18
c105 i9__carry_bar vss 42.7386e-18
c106 i9__net49 vss 123.595e-18
c107 i9__net51 vss 58.4059e-18
c108 i9__net50 vss 98.9679e-18
c109 i9__net52 vss 104.299e-18
c110 i7__net1 vss 83.3093e-18
c111 i7__carry_bar vss 42.7798e-18
c112 i7__net49 vss 124.38e-18
c113 i7__net51 vss 56.9149e-18
c114 i7__net50 vss 97.7831e-18
c115 i7__net52 vss 103.355e-18
c116 i10__net125 vss 117.881e-18
c117 i10__net122 vss 109.834e-18
c118 i10__net114 vss 80.6773e-18
c119 i10__net115 vss 86.871e-18
c120 i10__net124 vss 47.1088e-18
c121 i10__net116 vss 72.9089e-18
c122 i10__net118 vss 146.313e-18
c123 i10__net119 vss 144.087e-18
c124 i10__net121 vss 79.131e-18
c125 i10__net120 vss 80.373e-18
c126 i10__net117 vss 98.881e-18
c127 i10__net123 vss 75.7561e-18
c128 i2__net39 vss 73.3709e-18
c129 i2__net38 vss 99.1241e-18
c130 i2__net37 vss 77.5797e-18
c131 i2__net28 vss 96.9264e-18
c132 i2__net13 vss 78.3475e-18
c133 i2__net12 vss 98.3804e-18
c134 i2__net41 vss 79.5148e-18
c135 i2__net40 vss 96.8539e-18
c136 i2__net27 vss 76.0616e-18
c137 i2__net26 vss 98.3139e-18
c138 i2__net25 vss 77.5758e-18
c139 i2__net24 vss 95.7329e-18
c140 i2__net36 vss 79.0459e-18
c141 i2__net35 vss 104.986e-18
c142 i2__net34 vss 78.5737e-18
c143 i2__net33 vss 96.8322e-18
c144 i2__net2 vss 36.3036e-18
c145 i2__net4 vss 55.6198e-18
c146 i2__net3 vss 36.434e-18
c147 i2__rstb vss 16.2163e-18
c148 i2__net1 vss 36.295e-18
c149 i1__net39 vss 72.583e-18
c150 i1__net38 vss 99.5227e-18
c151 i1__net37 vss 77.458e-18
c152 i1__net28 vss 96.3985e-18
c153 i1__net13 vss 78.2e-18
c154 i1__net12 vss 101.422e-18
c155 i1__net41 vss 77.8307e-18
c156 i1__net40 vss 96.9101e-18
c157 i1__net27 vss 75.7663e-18
c158 i1__net26 vss 100.181e-18
c159 i1__net25 vss 77.983e-18
c160 i1__net24 vss 97.8828e-18
c161 i1__net36 vss 79.0384e-18
c162 i1__net35 vss 105.524e-18
c163 i1__net34 vss 81.7049e-18
c164 i1__net33 vss 95.7939e-18
c165 i1__net2 vss 37.5908e-18
c166 i1__net4 vss 55.6889e-18
c167 i1__net3 vss 36.3865e-18
c168 i1__rstb vss 17.4811e-18
c169 i1__net1 vss 36.9318e-18
c170 i0__net3 vss 31.7708e-18
c171 i0__net15 vss 94.4051e-18
c172 i0__net13 vss 98.9925e-18
c173 i0__net34 vss 97.5192e-18
c174 i0__net20 vss 89.9453e-18
c175 i0__net33 vss 86.8399e-18
c176 i0__net19 vss 101.853e-18
c177 i0__net17 vss 82.3945e-18
c178 i0__net16 vss 94.4845e-18
c179 i0__net6 vss 65.3608e-18
c180 i0__net4 vss 57.9456e-18
c181 i0__net2 vss 67.9047e-18
c182 i0__net1 vss 59.2294e-18
c183 n360__i12__net3 vss 338.944e-18
c184 n357__i12__net3 vss 291.96e-18
c185 n354__i12__net3 vss 285.122e-18
c186 n351__i12__net3 vss 285.021e-18
c187 n348__i12__net3 vss 285.209e-18
c188 n345__i12__net3 vss 284.983e-18
c189 n342__i12__net3 vss 285.063e-18
c190 n339__i12__net3 vss 285.369e-18
c191 n336__i12__net3 vss 285.063e-18
c192 n333__i12__net3 vss 284.983e-18
c193 n330__i12__net3 vss 285.209e-18
c194 n327__i12__net3 vss 284.983e-18
c195 n324__i12__net3 vss 285.063e-18
c196 n321__i12__net3 vss 285.369e-18
c197 n318__i12__net3 vss 285.063e-18
c198 n315__i12__net3 vss 284.983e-18
c199 n312__i12__net3 vss 285.209e-18
c200 n309__i12__net3 vss 284.983e-18
c201 n306__i12__net3 vss 285.063e-18
c202 n303__i12__net3 vss 285.369e-18
c203 n300__i12__net3 vss 285.063e-18
c204 n297__i12__net3 vss 285.021e-18
c205 n294__i12__net3 vss 285.483e-18
c206 n291__i12__net3 vss 285.305e-18
c207 n288__i12__net3 vss 285.261e-18
c208 n285__i12__net3 vss 285.724e-18
c209 n282__i12__net3 vss 285.408e-18
c210 n279__i12__net3 vss 285.217e-18
c211 n276__i12__net3 vss 285.507e-18
c212 n273__i12__net3 vss 285.235e-18
c213 n270__i12__net3 vss 285.261e-18
c214 n267__i12__net3 vss 285.724e-18
c215 n264__i12__net3 vss 285.408e-18
c216 n261__i12__net3 vss 285.217e-18
c217 n258__i12__net3 vss 285.507e-18
c218 n255__i12__net3 vss 285.235e-18
c219 n252__i12__net3 vss 285.261e-18
c220 n249__i12__net3 vss 285.724e-18
c221 n246__i12__net3 vss 285.408e-18
c222 n243__i12__net3 vss 285.217e-18
c223 n240__i12__net3 vss 285.507e-18
c224 n237__i12__net3 vss 285.235e-18
c225 n234__i12__net3 vss 285.261e-18
c226 n231__i12__net3 vss 285.724e-18
c227 n228__i12__net3 vss 285.708e-18
c228 n225__i12__net3 vss 285.444e-18
c229 n222__i12__net3 vss 285.163e-18
c230 n219__i12__net3 vss 284.878e-18
c231 n216__i12__net3 vss 284.754e-18
c232 n213__i12__net3 vss 285.009e-18
c233 n210__i12__net3 vss 285.392e-18
c234 n207__i12__net3 vss 285.246e-18
c235 n204__i12__net3 vss 285.094e-18
c236 n201__i12__net3 vss 285.427e-18
c237 n198__i12__net3 vss 285.286e-18
c238 n195__i12__net3 vss 285.5e-18
c239 n192__i12__net3 vss 286.418e-18
c240 n189__i12__net3 vss 286.244e-18
c241 n186__i12__net3 vss 285.509e-18
c242 n183__i12__net3 vss 285.532e-18
c243 n180__i12__net3 vss 285.217e-18
c244 n177__i12__net3 vss 285.009e-18
c245 n174__i12__net3 vss 285.392e-18
c246 n171__i12__net3 vss 285.246e-18
c247 n168__i12__net3 vss 285.094e-18
c248 n165__i12__net3 vss 285.298e-18
c249 n162__i12__net3 vss 285.067e-18
c250 n159__i12__net3 vss 285.096e-18
c251 n156__i12__net3 vss 285.447e-18
c252 n153__i12__net3 vss 285.03e-18
c253 n150__i12__net3 vss 285.107e-18
c254 n147__i12__net3 vss 285.569e-18
c255 n144__i12__net3 vss 285.239e-18
c256 n141__i12__net3 vss 285.393e-18
c257 n138__i12__net3 vss 285.567e-18
c258 n135__i12__net3 vss 284.951e-18
c259 n132__i12__net3 vss 285.107e-18
c260 n129__i12__net3 vss 285.569e-18
c261 n126__i12__net3 vss 285.239e-18
c262 n123__i12__net3 vss 285.38e-18
c263 n120__i12__net3 vss 285.438e-18
c264 n117__i12__net3 vss 284.911e-18
c265 n114__i12__net3 vss 285.063e-18
c266 n111__i12__net3 vss 285.369e-18
c267 n108__i12__net3 vss 285.063e-18
c268 n105__i12__net3 vss 284.983e-18
c269 n102__i12__net3 vss 285.209e-18
c270 n89__i12__net3 vss 284.983e-18
c271 n86__i12__net3 vss 285.063e-18
c272 n73__i12__net3 vss 285.369e-18
c273 n70__i12__net3 vss 285.063e-18
c274 n57__i12__net3 vss 284.954e-18
c275 n54__i12__net3 vss 284.974e-18
c276 n41__i12__net3 vss 284.723e-18
c277 n38__i12__net3 vss 285.048e-18
c278 n25__i12__net3 vss 289.317e-18
c279 n22__i12__net3 vss 311.573e-18
c280 n9__i12__net3 vss 285.3e-18
c281 n6__i12__net3 vss 288.189e-18
c282 n3__i12__net3 vss 320.532e-18
c283 n40__i12__net2 vss 394.031e-18
c284 n30__i12__net2 vss 320.897e-18
c285 n27__i12__net2 vss 319.182e-18
c286 n24__i12__net2 vss 287.65e-18
c287 n21__i12__net2 vss 287.741e-18
c288 n18__i12__net2 vss 287.648e-18
c289 n15__i12__net2 vss 287.788e-18
c290 n12__i12__net2 vss 287.782e-18
c291 n9__i12__net2 vss 287.454e-18
c292 n6__i12__net2 vss 291.186e-18
c293 n3__i12__net2 vss 341.023e-18
c294 n6__i12__net1 vss 231.685e-18
c295 n3__i12__net1 vss 244.32e-18
c296 n5__r_in vss 88.0435e-18
c297 n2__net5 vss 77.4681e-18
c298 n2__r_in vss 79.8125e-18
c299 n3__serial_out vss 28.7602e-18
c300 n25__clk vss 33.6522e-18
c301 n2__i14__net14 vss 56.8733e-18
c302 n24__i14__shift vss 36.9408e-18
c303 n21__clkb vss 34.0026e-18
c304 n17__i14__shift vss 27.889e-18
c305 n60__rst vss 44.8531e-18
c306 n16__i14__shift vss 31.0516e-18
c307 n21__clk vss 37.6973e-18
c308 n2__i14__net8 vss 56.7149e-18
c309 n9__i14__shift vss 24.8049e-18
c310 n17__clkb vss 36.041e-18
c311 n8__i14__shift vss 33.1483e-18
c312 n54__rst vss 44.5966e-18
c313 n17__clk vss 31.8417e-18
c314 n2__i14__net2 vss 57.0289e-18
c315 n13__clkb vss 36.3764e-18
c316 n48__rst vss 43.926e-18
c317 n17__clk2 vss 45.8702e-18
c318 n69__clk4 vss 48.1996e-18
c319 n5__i10__net116 vss 51.6293e-18
c320 n2__i10__net114 vss 54.51e-18
c321 n13__c0 vss 64.7514e-18
c322 n13__c1 vss 88.4827e-18
c323 n9__net12 vss 78.2053e-18
c324 n6__s1 vss 59.0219e-18
c325 n9__c0 vss 45.0192e-18
c326 n6__s0 vss 41.3987e-18
c327 n9__c1 vss 64.3971e-18
c328 n5__net12 vss 79.8231e-18
c329 n5__c1 vss 83.5332e-18
c330 n5__c0 vss 89.7951e-18
c331 n3__s1 vss 53.5111e-18
c332 n3__s0 vss 54.6708e-18
c333 n6__a1 vss 58.7425e-18
c334 n6__a3 vss 61.8268e-18
c335 n10__a0 vss 41.6591e-18
c336 n10__a2 vss 42.1367e-18
c337 n3__a1 vss 53.7892e-18
c338 n3__a3 vss 53.7781e-18
c339 n5__a0 vss 47.6566e-18
c340 n7__a0 vss 56.3936e-18
c341 n5__a2 vss 47.4875e-18
c342 n7__a2 vss 57.1515e-18
c343 n7__y1 vss 55.7091e-18
c344 n25__rst vss 46.5804e-18
c345 n21__rst vss 45.0732e-18
c346 n8__i1__rstb vss 28.2986e-18
c347 n8__i2__rstb vss 26.5514e-18
c348 n4__x1 vss 47.7079e-18
c349 n35__clk4b vss 34.7316e-18
c350 n33__clk4b vss 34.3356e-18
c351 n4__y3 vss 61.1432e-18
c352 n2__i1__net2 vss 56.5185e-18
c353 n2__i2__net2 vss 56.5442e-18
c354 n1__xin3 vss 58.245e-18
c355 n1__yin3 vss 58.4311e-18
c356 n32__clk4 vss 39.6375e-18
c357 n30__clk4 vss 40.886e-18
c358 n4__x3 vss 46.5564e-18
c359 n5__i1__rstb vss 29.3415e-18
c360 n5__i2__rstb vss 29.8506e-18
c361 n23__clk4b vss 32.9079e-18
c362 n21__clk4b vss 32.6199e-18
c363 n1__xin2 vss 57.9267e-18
c364 n1__yin2 vss 57.6196e-18
c365 n24__clk4 vss 33.9736e-18
c366 n22__clk4 vss 33.6993e-18
c367 n15__clk4b vss 36.2894e-18
c368 n13__clk4b vss 34.8774e-18
c369 n2__i1__net3 vss 55.8168e-18
c370 n2__i2__net3 vss 55.8136e-18
c371 n1__xin1 vss 57.7895e-18
c372 n1__yin1 vss 57.8119e-18
c373 n16__clk4 vss 41.0487e-18
c374 n14__clk4 vss 41.0245e-18
c375 n3__i1__rstb vss 25.7906e-18
c376 n3__i2__rstb vss 25.7207e-18
c377 n4__y0 vss 56.8173e-18
c378 n4__y2 vss 58.6132e-18
c379 n4__x0 vss 47.5324e-18
c380 n7__clk4b vss 32.7956e-18
c381 n5__clk4b vss 31.8709e-18
c382 n4__x2 vss 47.0564e-18
c383 n2__i1__net1 vss 56.2034e-18
c384 n2__i2__net1 vss 55.863e-18
c385 n1__xin0 vss 57.5731e-18
c386 n1__yin0 vss 57.7474e-18
c387 n8__clk4 vss 30.4394e-18
c388 n6__clk4 vss 33.1636e-18
c389 n4__i0__net4 vss 30.0673e-18
c390 n6__i0__net1 vss 33.5613e-18
c391 n2__i0__net6 vss 56.9346e-18
c392 n6__clk2 vss 32.5746e-18
c393 n3__clkb vss 32.4311e-18
c394 n2__i0__net2 vss 57.3362e-18
c395 n3__clk vss 46.0376e-18
c396 n2__clk vss 36.147e-18
c397 n359__i12__net3 vss 204.238e-18
c398 n356__i12__net3 vss 166.952e-18
c399 n353__i12__net3 vss 164.305e-18
c400 n350__i12__net3 vss 164.123e-18
c401 n347__i12__net3 vss 164.17e-18
c402 n344__i12__net3 vss 163.944e-18
c403 n341__i12__net3 vss 164.024e-18
c404 n338__i12__net3 vss 164.329e-18
c405 n335__i12__net3 vss 164.024e-18
c406 n332__i12__net3 vss 163.944e-18
c407 n329__i12__net3 vss 164.17e-18
c408 n326__i12__net3 vss 163.944e-18
c409 n323__i12__net3 vss 164.024e-18
c410 n320__i12__net3 vss 164.329e-18
c411 n317__i12__net3 vss 164.024e-18
c412 n314__i12__net3 vss 163.944e-18
c413 n311__i12__net3 vss 164.17e-18
c414 n308__i12__net3 vss 163.944e-18
c415 n305__i12__net3 vss 164.024e-18
c416 n302__i12__net3 vss 164.329e-18
c417 n299__i12__net3 vss 164.024e-18
c418 n296__i12__net3 vss 163.982e-18
c419 n293__i12__net3 vss 164.444e-18
c420 n290__i12__net3 vss 164.266e-18
c421 n287__i12__net3 vss 164.222e-18
c422 n284__i12__net3 vss 164.685e-18
c423 n281__i12__net3 vss 164.369e-18
c424 n278__i12__net3 vss 164.177e-18
c425 n275__i12__net3 vss 164.468e-18
c426 n272__i12__net3 vss 164.196e-18
c427 n269__i12__net3 vss 164.222e-18
c428 n266__i12__net3 vss 164.685e-18
c429 n263__i12__net3 vss 164.369e-18
c430 n260__i12__net3 vss 164.177e-18
c431 n257__i12__net3 vss 164.468e-18
c432 n254__i12__net3 vss 164.196e-18
c433 n251__i12__net3 vss 164.222e-18
c434 n248__i12__net3 vss 164.685e-18
c435 n245__i12__net3 vss 164.369e-18
c436 n242__i12__net3 vss 164.177e-18
c437 n239__i12__net3 vss 164.468e-18
c438 n236__i12__net3 vss 164.196e-18
c439 n233__i12__net3 vss 164.222e-18
c440 n230__i12__net3 vss 164.685e-18
c441 n227__i12__net3 vss 164.668e-18
c442 n224__i12__net3 vss 164.404e-18
c443 n221__i12__net3 vss 164.123e-18
c444 n218__i12__net3 vss 163.839e-18
c445 n215__i12__net3 vss 163.715e-18
c446 n212__i12__net3 vss 163.97e-18
c447 n209__i12__net3 vss 164.353e-18
c448 n206__i12__net3 vss 164.207e-18
c449 n203__i12__net3 vss 164.055e-18
c450 n200__i12__net3 vss 164.378e-18
c451 n197__i12__net3 vss 164.216e-18
c452 n194__i12__net3 vss 164.339e-18
c453 n191__i12__net3 vss 165.99e-18
c454 n188__i12__net3 vss 166.427e-18
c455 n185__i12__net3 vss 164.47e-18
c456 n182__i12__net3 vss 164.493e-18
c457 n179__i12__net3 vss 164.177e-18
c458 n176__i12__net3 vss 163.97e-18
c459 n173__i12__net3 vss 164.353e-18
c460 n170__i12__net3 vss 164.207e-18
c461 n167__i12__net3 vss 164.055e-18
c462 n164__i12__net3 vss 164.259e-18
c463 n161__i12__net3 vss 164.028e-18
c464 n158__i12__net3 vss 164.056e-18
c465 n155__i12__net3 vss 164.408e-18
c466 n152__i12__net3 vss 163.99e-18
c467 n149__i12__net3 vss 164.068e-18
c468 n146__i12__net3 vss 164.53e-18
c469 n143__i12__net3 vss 164.2e-18
c470 n140__i12__net3 vss 164.354e-18
c471 n137__i12__net3 vss 164.528e-18
c472 n134__i12__net3 vss 163.912e-18
c473 n131__i12__net3 vss 164.068e-18
c474 n128__i12__net3 vss 164.53e-18
c475 n125__i12__net3 vss 164.2e-18
c476 n122__i12__net3 vss 164.341e-18
c477 n119__i12__net3 vss 164.399e-18
c478 n116__i12__net3 vss 163.872e-18
c479 n113__i12__net3 vss 164.024e-18
c480 n110__i12__net3 vss 164.329e-18
c481 n107__i12__net3 vss 164.024e-18
c482 n104__i12__net3 vss 163.944e-18
c483 n101__i12__net3 vss 164.17e-18
c484 n88__i12__net3 vss 163.944e-18
c485 n85__i12__net3 vss 164.024e-18
c486 n72__i12__net3 vss 164.329e-18
c487 n69__i12__net3 vss 164.024e-18
c488 n56__i12__net3 vss 163.915e-18
c489 n53__i12__net3 vss 163.935e-18
c490 n40__i12__net3 vss 163.681e-18
c491 n37__i12__net3 vss 164.008e-18
c492 n24__i12__net3 vss 166.442e-18
c493 n21__i12__net3 vss 178.948e-18
c494 n8__i12__net3 vss 164.259e-18
c495 n5__i12__net3 vss 165.46e-18
c496 n2__i12__net3 vss 181.57e-18
c497 n39__i12__net2 vss 202.748e-18
c498 n29__i12__net2 vss 204.623e-18
c499 n26__i12__net2 vss 164.318e-18
c500 n23__i12__net2 vss 164.003e-18
c501 n20__i12__net2 vss 163.951e-18
c502 n17__i12__net2 vss 163.859e-18
c503 n14__i12__net2 vss 163.998e-18
c504 n11__i12__net2 vss 163.992e-18
c505 n8__i12__net2 vss 163.664e-18
c506 n5__i12__net2 vss 164.883e-18
c507 n2__i12__net2 vss 191.905e-18
c508 n5__i12__net1 vss 142.978e-18
c509 n2__i12__net1 vss 150.177e-18
c510 n4__r_in vss 57.4537e-18
c511 n2__i11__net1 vss 159.108e-18
c512 n2__serial_out vss 197.514e-18
c513 n5__serial_out vss 34.9134e-18
c514 n22__clkb vss 26.5979e-18
c515 n3__i14__net14 vss 61.2831e-18
c516 n3__i14__i2__net1 vss 28.3214e-18
c517 n3__i14__i5__net5 vss 59.7845e-18
c518 n21__i14__shift vss 32.1414e-18
c519 n24__clk vss 27.3442e-18
c520 n20__i14__shift vss 20.5033e-18
c521 n62__rst vss 18.6287e-18
c522 n59__rst vss 20.3045e-18
c523 n3__i14__i1__net1 vss 30.2408e-18
c524 n13__i14__shift vss 32.0599e-18
c525 n18__clkb vss 26.2022e-18
c526 n3__i14__net8 vss 63.6258e-18
c527 n12__i14__shift vss 17.5783e-18
c528 n3__i14__i4__net5 vss 60.1338e-18
c529 n20__clk vss 27.9021e-18
c530 n3__i14__i0__net1 vss 29.8247e-18
c531 n5__i14__shift vss 32.334e-18
c532 n56__rst vss 19.1845e-18
c533 n53__rst vss 18.4169e-18
c534 n4__i14__shift vss 17.1657e-18
c535 n14__clkb vss 25.9787e-18
c536 n3__i14__net2 vss 63.5689e-18
c537 n3__i14__i3__net5 vss 59.9182e-18
c538 n16__clk vss 27.8586e-18
c539 n4__i14__i7__net1 vss 26.3308e-18
c540 n50__rst vss 18.849e-18
c541 n47__rst vss 16.541e-18
c542 n19__clk2 vss 31.2121e-18
c543 n71__clk4 vss 31.348e-18
c544 n8__i10__net116 vss 25.0111e-18
c545 n3__i10__net114 vss 45.7466e-18
c546 n16__c0 vss 67.4261e-18
c547 n16__c1 vss 63.0595e-18
c548 n12__net12 vss 46.3932e-18
c549 n8__s1 vss 77.9397e-18
c550 n12__c0 vss 54.8013e-18
c551 n8__s0 vss 92.8727e-18
c552 n12__c1 vss 57.1308e-18
c553 n8__net12 vss 45.3489e-18
c554 n3__i9__carry_bar vss 59.5852e-18
c555 n4__i10__net116 vss 29.6302e-18
c556 n3__i9__net51 vss 48.4389e-18
c557 n8__c1 vss 63.8926e-18
c558 n8__c0 vss 82.2925e-18
c559 n4__net12 vss 46.9021e-18
c560 n4__s1 vss 46.2136e-18
c561 n5__s1 vss 33.1864e-18
c562 n4__s0 vss 42.1562e-18
c563 n5__s0 vss 34.703e-18
c564 n4__c1 vss 49.064e-18
c565 n4__c0 vss 52.9032e-18
c566 n8__a1 vss 71.7372e-18
c567 n8__a3 vss 79.9402e-18
c568 n12__a0 vss 96.9872e-18
c569 n12__a2 vss 96.9712e-18
c570 n3__i7__carry_bar vss 58.7623e-18
c571 n3__i8__carry_bar vss 63.0812e-18
c572 n3__i7__net51 vss 48.4565e-18
c573 n3__i8__net51 vss 48.268e-18
c574 n4__a1 vss 46.6277e-18
c575 n5__a1 vss 38.405e-18
c576 n4__a3 vss 46.667e-18
c577 n5__a3 vss 38.086e-18
c578 n8__a0 vss 42.6878e-18
c579 n9__a0 vss 35.2084e-18
c580 n8__a2 vss 41.2236e-18
c581 n9__a2 vss 34.9162e-18
c582 n10__y1 vss 32.7908e-18
c583 n28__rst vss 19.7791e-18
c584 n24__rst vss 16.7774e-18
c585 n3__i4__abar vss 71.9529e-18
c586 n15__rst vss 15.0417e-18
c587 n13__rst vss 14.5176e-18
c588 n3__i4__bbar vss 64.2571e-18
c589 n7__x1 vss 45.4334e-18
c590 n39__clk4 vss 25.5784e-18
c591 n37__clk4 vss 26.263e-18
c592 n7__y3 vss 29.1145e-18
c593 n3__i1__net2 vss 58.2073e-18
c594 n3__i2__net2 vss 58.626e-18
c595 n3__i6__abar vss 70.5303e-18
c596 n3__y1 vss 30.871e-18
c597 n3__xin3 vss 62.457e-18
c598 n3__yin3 vss 58.736e-18
c599 n3__i6__bbar vss 65.9492e-18
c600 n3__x1 vss 40.1056e-18
c601 n28__clk4b vss 24.3822e-18
c602 n26__clk4b vss 23.4217e-18
c603 n7__x3 vss 44.191e-18
c604 n11__rst vss 29.8292e-18
c605 n9__rst vss 26.6641e-18
c606 n3__y3 vss 31.7254e-18
c607 n27__clk4 vss 38.5217e-18
c608 n25__clk4 vss 37.721e-18
c609 n3__x3 vss 45.8051e-18
c610 n2__i1__net4 vss 63.8846e-18
c611 n2__i2__net4 vss 64.5426e-18
c612 n3__xin2 vss 62.2189e-18
c613 n3__yin2 vss 59.2785e-18
c614 n20__clk4b vss 22.9037e-18
c615 n18__clk4b vss 23.3525e-18
c616 n19__clk4 vss 25.1425e-18
c617 n17__clk4 vss 24.7336e-18
c618 n3__i1__net3 vss 59.8441e-18
c619 n3__i2__net3 vss 58.3222e-18
c620 n3__xin1 vss 61.1173e-18
c621 n3__yin1 vss 59.1548e-18
c622 n12__clk4b vss 20.9713e-18
c623 n10__clk4b vss 21.9477e-18
c624 n7__y0 vss 30.4287e-18
c625 n7__y2 vss 30.8056e-18
c626 n3__i3__abar vss 71.9686e-18
c627 n8__rst vss 14.8742e-18
c628 n6__rst vss 14.3413e-18
c629 n3__i5__abar vss 72.8103e-18
c630 n3__i3__bbar vss 64.3167e-18
c631 n3__rst vss 19.8992e-18
c632 n1__rst vss 19.4553e-18
c633 n3__i5__bbar vss 64.8701e-18
c634 n7__x0 vss 45.5709e-18
c635 n11__clk4 vss 38.2261e-18
c636 n9__clk4 vss 38.1178e-18
c637 n7__x2 vss 45.7047e-18
c638 n3__i1__net1 vss 59.2285e-18
c639 n3__i2__net1 vss 60.6948e-18
c640 n3__y0 vss 31.1719e-18
c641 n3__xin0 vss 60.6653e-18
c642 n3__yin0 vss 61.7066e-18
c643 n3__y2 vss 31.934e-18
c644 n3__x0 vss 40.5368e-18
c645 n4__clk4b vss 23.4895e-18
c646 n2__clk4b vss 27.1708e-18
c647 n3__x2 vss 41.3299e-18
c648 n4__clk4 vss 22.1988e-18
c649 n7__i0__net4 vss 21.637e-18
c650 n4__i0__net3 vss 20.2671e-18
c651 n7__clk2 vss 26.5919e-18
c652 n3__i0__net6 vss 59.1694e-18
c653 n3__i0__net4 vss 63.4601e-18
c654 n5__i0__net1 vss 23.1477e-18
c655 n4__clk2 vss 17.825e-18
c656 n7__clk vss 24.8482e-18
c657 n3__i0__net2 vss 61.2087e-18
c658 n6__clk vss 32.7612e-18
c659 n3__i0__net1 vss 63.7335e-18
c660 n2__clkb vss 25.0864e-18
c661 n358__i12__net3 vss 58.5487e-18
c662 n355__i12__net3 vss 43.4935e-18
c663 n352__i12__net3 vss 43.014e-18
c664 n349__i12__net3 vss 42.7716e-18
c665 n346__i12__net3 vss 42.6442e-18
c666 n343__i12__net3 vss 42.6063e-18
c667 n340__i12__net3 vss 42.5323e-18
c668 n337__i12__net3 vss 42.5489e-18
c669 n334__i12__net3 vss 42.5881e-18
c670 n331__i12__net3 vss 42.4944e-18
c671 n328__i12__net3 vss 42.6442e-18
c672 n325__i12__net3 vss 42.6063e-18
c673 n322__i12__net3 vss 42.5323e-18
c674 n319__i12__net3 vss 42.5489e-18
c675 n316__i12__net3 vss 42.5881e-18
c676 n313__i12__net3 vss 42.4944e-18
c677 n310__i12__net3 vss 42.6442e-18
c678 n307__i12__net3 vss 42.6063e-18
c679 n304__i12__net3 vss 42.5323e-18
c680 n301__i12__net3 vss 42.5489e-18
c681 n298__i12__net3 vss 42.5881e-18
c682 n295__i12__net3 vss 42.4944e-18
c683 n292__i12__net3 vss 42.6442e-18
c684 n289__i12__net3 vss 42.4384e-18
c685 n286__i12__net3 vss 42.8446e-18
c686 n283__i12__net3 vss 43.5019e-18
c687 n280__i12__net3 vss 42.7413e-18
c688 n277__i12__net3 vss 43.5607e-18
c689 n274__i12__net3 vss 42.7972e-18
c690 n271__i12__net3 vss 42.4384e-18
c691 n268__i12__net3 vss 42.8446e-18
c692 n265__i12__net3 vss 43.5019e-18
c693 n262__i12__net3 vss 42.7413e-18
c694 n259__i12__net3 vss 43.5607e-18
c695 n256__i12__net3 vss 42.7972e-18
c696 n253__i12__net3 vss 42.4384e-18
c697 n250__i12__net3 vss 42.8446e-18
c698 n247__i12__net3 vss 43.5019e-18
c699 n244__i12__net3 vss 42.7413e-18
c700 n241__i12__net3 vss 43.5607e-18
c701 n238__i12__net3 vss 42.7972e-18
c702 n235__i12__net3 vss 42.4384e-18
c703 n232__i12__net3 vss 42.8446e-18
c704 n229__i12__net3 vss 43.5019e-18
c705 n226__i12__net3 vss 42.7413e-18
c706 n223__i12__net3 vss 43.5607e-18
c707 n220__i12__net3 vss 42.7972e-18
c708 n217__i12__net3 vss 42.6049e-18
c709 n214__i12__net3 vss 42.5321e-18
c710 n211__i12__net3 vss 42.5504e-18
c711 n208__i12__net3 vss 42.5882e-18
c712 n205__i12__net3 vss 42.8067e-18
c713 n202__i12__net3 vss 42.4763e-18
c714 n199__i12__net3 vss 42.6049e-18
c715 n196__i12__net3 vss 42.5321e-18
c716 n193__i12__net3 vss 42.5504e-18
c717 n190__i12__net3 vss 42.5882e-18
c718 n187__i12__net3 vss 42.8067e-18
c719 n184__i12__net3 vss 42.4763e-18
c720 n181__i12__net3 vss 42.6049e-18
c721 n178__i12__net3 vss 42.5321e-18
c722 n175__i12__net3 vss 42.5504e-18
c723 n172__i12__net3 vss 42.5882e-18
c724 n169__i12__net3 vss 42.8067e-18
c725 n166__i12__net3 vss 42.4763e-18
c726 n163__i12__net3 vss 42.6049e-18
c727 n160__i12__net3 vss 42.5321e-18
c728 n157__i12__net3 vss 42.5504e-18
c729 n154__i12__net3 vss 42.5882e-18
c730 n151__i12__net3 vss 42.4944e-18
c731 n148__i12__net3 vss 42.6442e-18
c732 n145__i12__net3 vss 42.437e-18
c733 n142__i12__net3 vss 42.8434e-18
c734 n139__i12__net3 vss 43.512e-18
c735 n136__i12__net3 vss 42.7413e-18
c736 n133__i12__net3 vss 42.4944e-18
c737 n130__i12__net3 vss 42.6442e-18
c738 n127__i12__net3 vss 42.437e-18
c739 n124__i12__net3 vss 42.8434e-18
c740 n121__i12__net3 vss 43.512e-18
c741 n118__i12__net3 vss 42.7413e-18
c742 n115__i12__net3 vss 42.6063e-18
c743 n112__i12__net3 vss 42.5323e-18
c744 n109__i12__net3 vss 42.5489e-18
c745 n106__i12__net3 vss 42.5881e-18
c746 n103__i12__net3 vss 42.4944e-18
c747 n100__i12__net3 vss 42.6442e-18
c748 n87__i12__net3 vss 42.6063e-18
c749 n84__i12__net3 vss 42.5323e-18
c750 n71__i12__net3 vss 42.5489e-18
c751 n68__i12__net3 vss 42.5881e-18
c752 n55__i12__net3 vss 42.4944e-18
c753 n52__i12__net3 vss 42.6442e-18
c754 n39__i12__net3 vss 42.5504e-18
c755 n36__i12__net3 vss 42.5882e-18
c756 n23__i12__net3 vss 42.8067e-18
c757 n20__i12__net3 vss 42.4763e-18
c758 n7__i12__net3 vss 42.6049e-18
c759 n4__i12__net3 vss 42.1955e-18
c760 n38__i12__net2 vss 57.352e-18
c761 n28__i12__net2 vss 42.7368e-18
c762 n25__i12__net2 vss 42.0904e-18
c763 n22__i12__net2 vss 42.6905e-18
c764 n19__i12__net2 vss 41.7866e-18
c765 n16__i12__net2 vss 42.2293e-18
c766 n13__i12__net2 vss 41.7803e-18
c767 n10__i12__net2 vss 42.1049e-18
c768 n7__i12__net2 vss 41.7082e-18
c769 n4__i12__net2 vss 41.8126e-18
c770 n4__i12__net1 vss 58.6196e-18
c771 n3__r_in vss 165.925e-18
c772 n4__serial_out vss 78.3174e-18
c773 n23__clkb vss 98.8304e-18
c774 n26__clk vss 44.6935e-18
c775 n23__i14__shift vss 28.9217e-18
c776 n4__i14__i2__net1 vss 93.2412e-18
c777 n2__i14__i5__net5 vss 40.3216e-18
c778 n22__i14__shift vss 20.9221e-18
c779 n2__i14__i2__net1 vss 28.3287e-18
c780 n20__clkb vss 116.461e-18
c781 n23__clk vss 38.3564e-18
c782 n61__rst vss 53.9148e-18
c783 n19__i14__shift vss 11.5857e-18
c784 n2__i14__i5__rstb vss 86.8324e-18
c785 n57__rst vss 28.6773e-18
c786 n15__i14__shift vss 23.8809e-18
c787 n4__i14__i1__net1 vss 106.713e-18
c788 n14__i14__shift vss 19.2701e-18
c789 n2__i14__i1__net1 vss 26.8621e-18
c790 n19__clkb vss 102.128e-18
c791 n22__clk vss 45.362e-18
c792 n11__i14__shift vss 12.2137e-18
c793 n2__i14__i4__net5 vss 38.2525e-18
c794 n16__clkb vss 117.041e-18
c795 n19__clk vss 38.6597e-18
c796 n7__i14__shift vss 23.5827e-18
c797 n4__i14__i0__net1 vss 110.051e-18
c798 n55__rst vss 53.4575e-18
c799 n6__i14__shift vss 19.9781e-18
c800 n2__i14__i0__net1 vss 25.9916e-18
c801 n2__i14__i4__rstb vss 87.2426e-18
c802 n51__rst vss 128.355e-18
c803 n3__i14__shift vss 10.1142e-18
c804 n15__clkb vss 102.465e-18
c805 n18__clk vss 44.7902e-18
c806 n2__i14__i3__net5 vss 37.0721e-18
c807 n12__clkb vss 114.063e-18
c808 n15__clk vss 39.0519e-18
c809 n49__rst vss 51.7429e-18
c810 n3__i14__i7__net1 vss 23.5039e-18
c811 n2__i14__i3__rstb vss 84.5389e-18
c812 n45__rst vss 31.0407e-18
c813 n18__clk2 vss 36.1485e-18
c814 n70__clk4 vss 36.7156e-18
c815 n7__i10__net116 vss 47.2782e-18
c816 n6__i10__net114 vss 48.2959e-18
c817 n15__c0 vss 106.18e-18
c818 n15__c1 vss 143.571e-18
c819 n11__net12 vss 120.186e-18
c820 n7__s1 vss 94.7818e-18
c821 n11__c0 vss 237.47e-18
c822 n7__s0 vss 94.0353e-18
c823 n11__c1 vss 275.398e-18
c824 n7__net12 vss 276.379e-18
c825 n2__i9__carry_bar vss 109.437e-18
c826 n3__i10__net116 vss 13.1455e-18
c827 n2__i9__net51 vss 56.1302e-18
c828 n7__c1 vss 279.426e-18
c829 n7__c0 vss 239.654e-18
c830 n2__s1 vss 34.2566e-18
c831 n3__net12 vss 289.468e-18
c832 n2__s0 vss 33.4688e-18
c833 n3__c1 vss 191.361e-18
c834 n3__c0 vss 379.427e-18
c835 n7__a1 vss 82.2787e-18
c836 n7__a3 vss 94.4498e-18
c837 n11__a0 vss 98.226e-18
c838 n11__a2 vss 99.9567e-18
c839 n2__i7__carry_bar vss 110.595e-18
c840 n2__i8__carry_bar vss 109.678e-18
c841 n2__i7__net51 vss 56.6688e-18
c842 n2__i8__net51 vss 100.766e-18
c843 n2__a1 vss 35.4308e-18
c844 n2__a3 vss 34.6503e-18
c845 n6__a0 vss 34.5492e-18
c846 n6__a2 vss 34.2673e-18
c847 n9__y1 vss 45.9874e-18
c848 n27__rst vss 83.4209e-18
c849 n23__rst vss 86.9205e-18
c850 n7__i1__rstb vss 36.2329e-18
c851 n7__i2__rstb vss 36.7319e-18
c852 n2__i4__abar vss 310.823e-18
c853 n16__rst vss 21.0867e-18
c854 n14__rst vss 20.65e-18
c855 n2__i4__bbar vss 176.332e-18
c856 n6__x1 vss 67.2902e-18
c857 n40__clk4 vss 39.0842e-18
c858 n38__clk4 vss 40.2024e-18
c859 n36__clk4b vss 116.358e-18
c860 n34__clk4b vss 117.916e-18
c861 n6__y3 vss 40.5402e-18
c862 n2__i6__abar vss 312.428e-18
c863 n2__y1 vss 33.5483e-18
c864 n2__xin3 vss 74.0933e-18
c865 n2__yin3 vss 35.2616e-18
c866 n2__i6__bbar vss 173.413e-18
c867 n31__clk4 vss 46.8295e-18
c868 n27__clk4b vss 92.7055e-18
c869 n29__clk4 vss 46.4717e-18
c870 n25__clk4b vss 92.6574e-18
c871 n2__x1 vss 36.2263e-18
c872 n6__x3 vss 71.1825e-18
c873 n6__i1__rstb vss 22.595e-18
c874 n6__i2__rstb vss 23.9848e-18
c875 n2__y3 vss 33.4707e-18
c876 n12__rst vss 33.5862e-18
c877 n10__rst vss 33.5125e-18
c878 n24__clk4b vss 121.776e-18
c879 n28__clk4 vss 94.0186e-18
c880 n2__x3 vss 37.1917e-18
c881 n22__clk4b vss 122.068e-18
c882 n26__clk4 vss 46.4741e-18
c883 n3__i1__net4 vss 69.9827e-18
c884 n3__i2__net4 vss 36.6797e-18
c885 n2__xin2 vss 83.8022e-18
c886 n2__yin2 vss 91.5499e-18
c887 n23__clk4 vss 42.5675e-18
c888 n19__clk4b vss 95.6312e-18
c889 n21__clk4 vss 42.0045e-18
c890 n17__clk4b vss 95.3481e-18
c891 n20__clk4 vss 38.262e-18
c892 n18__clk4 vss 38.863e-18
c893 n16__clk4b vss 113.612e-18
c894 n14__clk4b vss 115.02e-18
c895 n2__xin1 vss 82.0902e-18
c896 n2__yin1 vss 35.3982e-18
c897 n15__clk4 vss 47.8353e-18
c898 n11__clk4b vss 92.5429e-18
c899 n13__clk4 vss 47.3713e-18
c900 n9__clk4b vss 92.6171e-18
c901 n4__i1__rstb vss 20.2174e-18
c902 n4__i2__rstb vss 20.6143e-18
c903 n2__i1__rstb vss 50.765e-18
c904 n2__i2__rstb vss 49.5075e-18
c905 n6__y0 vss 69.4244e-18
c906 n6__y2 vss 38.4681e-18
c907 n7__rst vss 22.125e-18
c908 n5__rst vss 20.4303e-18
c909 n2__i3__abar vss 311.16e-18
c910 n2__i5__abar vss 312.769e-18
c911 n2__i3__bbar vss 175.481e-18
c912 n4__rst vss 29.3663e-18
c913 n2__rst vss 29.1016e-18
c914 n2__i5__bbar vss 173.491e-18
c915 n6__x0 vss 38.3662e-18
c916 n12__clk4 vss 40.2276e-18
c917 n10__clk4 vss 41.5525e-18
c918 n8__clk4b vss 113.974e-18
c919 n6__clk4b vss 114.639e-18
c920 n6__x2 vss 39.0665e-18
c921 n2__y0 vss 33.359e-18
c922 n2__xin0 vss 76.2885e-18
c923 n2__yin0 vss 32.9736e-18
c924 n2__y2 vss 34.694e-18
c925 n7__clk4 vss 40.6111e-18
c926 n3__clk4b vss 104.501e-18
c927 n5__clk4 vss 43.1314e-18
c928 n2__x0 vss 35.9763e-18
c929 n2__x2 vss 36.1372e-18
c930 n3__clk4 vss 69.0464e-18
c931 n6__i0__net4 vss 73.5829e-18
c932 n3__i0__net3 vss 77.4653e-18
c933 n8__clk2 vss 38.7869e-18
c934 n7__i0__net1 vss 153.493e-18
c935 n2__i0__net4 vss 87.0751e-18
c936 n5__clk2 vss 39.8938e-18
c937 n4__i0__net1 vss 38.2247e-18
c938 n3__clk2 vss 71.2034e-18
c939 n8__clk vss 37.7137e-18
c940 n4__clkb vss 149.445e-18
c941 n5__clk vss 106.006e-18
c942 n2__i0__net1 vss 86.6936e-18
c943 n1__clk vss 42.9788e-18
c944 n282__vdd vss 745.983e-18
c945 n314__vddio vss 41.0685e-18
c946 n247__vdd vss 567.876e-18
c947 n246__vdd vss 402.808e-18
c948 n184__vdd vss 361.711e-18
c949 n95__vdd vss 349.763e-18
c950 n52__vdd vss 409.932e-18
c951 n13__vdd vss 191.415e-18
c952 n311__vddio vss 1.13883e-18
c953 n281__vdd vss 157.034e-18
c954 n310__vddio vss 76.7036e-18
c955 n245__vdd vss 70.666e-18
c956 n243__vdd vss 101.654e-18
c957 n244__vdd vss 279.623e-18
c958 n183__vdd vss 111.806e-18
c959 n94__vdd vss 100.913e-18
c960 n92__vdd vss 58.3244e-18
c961 n89__vdd vss 130.609e-18
c962 n46__vdd vss 70.8965e-18
c963 n49__vdd vss 59.2545e-18
c964 n50__vdd vss 96.6335e-18
c965 n45__vdd vss 5.7639e-18
c966 n12__vdd vss 30.1446e-18
c967 n309__vddio vss 2.39802e-18
c968 n280__vdd vss 13.5163e-18
c969 n242__vdd vss 358.04e-21
c970 n226__vdd vss 2.45846e-18
c971 n227__vdd vss 3.37337e-18
c972 n143__vdd vss 6.22933e-18
c973 n140__vdd vss 314.084e-18
c974 n11__vdd vss 12.059e-18
c975 n279__vdd vss 6.25131e-18
c976 n306__vddio vss 1.45471e-18
c977 n17__r0 vss 253.407e-18
c978 n9__r0 vss 320.942e-18
c979 n225__vdd vss 6.06233e-18
c980 n142__vdd vss 7.40785e-18
c981 n141__vdd vss 4.31305e-18
c982 n88__vdd vss 25.9505e-18
c983 n87__vdd vss 7.46299e-18
c984 n41__vdd vss 11.162e-18
c985 n42__vdd vss 8.3036e-18
c986 n43__vdd vss 1.61457e-18
c987 n40__vdd vss 7.66171e-18
c988 n9__vdd vss 6.54168e-18
c989 n240__vdd vss 3.14081e-18
c990 n65__rst vss 317.343e-18
c991 n205__vdd vss 1.39648e-18
c992 n206__vdd vss 5.23255e-18
c993 n44__rst vss 47.0404e-18
c994 n33__rst vss 254.13e-18
c995 n85__vdd vss 11.0841e-18
c996 n83__vdd vss 14.2322e-18
c997 n37__vdd vss 1.67926e-18
c998 n38__vdd vss 8.78276e-18
c999 n39__vdd vss 5.73053e-18
c1000 n36__vdd vss 11.8527e-18
c1001 n277__vdd vss 7.6887e-18
c1002 n15__r0 vss 678.897e-21
c1003 n12__r1 vss 131.991e-18
c1004 n34__clk vss 141.896e-18
c1005 n239__vdd vss 21.8087e-18
c1006 n66__rst vss 29.929e-18
c1007 n7__r1 vss 179.468e-18
c1008 n7__r0 vss 70.3784e-18
c1009 n189__vdd vss 1.33455e-18
c1010 n190__vdd vss 11.1607e-18
c1011 n147__vdd vss 15.3941e-18
c1012 n144__vdd vss 14.5296e-18
c1013 n34__rst vss 13.4625e-18
c1014 n32__rst vss 6.91659e-18
c1015 n82__vdd vss 9.15135e-18
c1016 n80__vdd vss 85.9645e-18
c1017 n34__vdd vss 63.7733e-18
c1018 n35__vdd vss 45.7416e-18
c1019 n3__vdd vss 5.14418e-18
c1020 n9__clk vss 273.833e-18
c1021 n269__vdd vss 10.5163e-18
c1022 n13__serial_out vss 79.0089e-18
c1023 n14__r0 vss 3.66954e-18
c1024 n7__i14__net14 vss 96.2694e-18
c1025 n9__i14__net14 vss 74.4956e-18
c1026 n10__i14__net15 vss 206.745e-18
c1027 n11__serial_out vss 28.2854e-18
c1028 n11__r1 vss 48.0849e-18
c1029 n71__rst vss 129.718e-18
c1030 n8__i14__net8 vss 115.898e-18
c1031 n9__i14__net8 vss 100.723e-18
c1032 n10__i14__net9 vss 215.22e-18
c1033 n6__i14__net15 vss 226.029e-18
c1034 n9__r2 vss 165.987e-18
c1035 n4__i14__net2 vss 118.603e-18
c1036 n5__i14__net2 vss 90.9227e-18
c1037 n69__rst vss 56.3133e-18
c1038 n6__i14__net9 vss 207.501e-18
c1039 n28__clk vss 19.1671e-18
c1040 n237__vdd vss 79.255e-18
c1041 n238__vdd vss 71.923e-18
c1042 n64__rst vss 39.3541e-18
c1043 n22__clk2 vss 1.08608e-15
c1044 n74__clk4 vss 986.022e-18
c1045 n5__r2 vss 212.453e-18
c1046 n185__vdd vss 4.8549e-18
c1047 n188__vdd vss 19.3478e-18
c1048 n6__r0 vss 75.8881e-18
c1049 n15__s1 vss 397.029e-18
c1050 n14__s1 vss 230.32e-18
c1051 n35__rst vss 19.3151e-18
c1052 n31__rst vss 41.6301e-18
c1053 n14__x3 vss 253.927e-18
c1054 n15__y3 vss 237.967e-18
c1055 n21__y1 vss 334.692e-18
c1056 n77__vdd vss 32.4047e-18
c1057 n69__vdd vss 21.6329e-18
c1058 n24__x1 vss 325.999e-18
c1059 n13__y3 vss 319.775e-18
c1060 n18__x2 vss 284.668e-18
c1061 n18__y2 vss 365.94e-18
c1062 n13__x3 vss 229.981e-18
c1063 n18__x1 vss 128.718e-18
c1064 n18__y1 vss 143.443e-18
c1065 n12__x1 vss 223.957e-18
c1066 n12__y1 vss 199.688e-18
c1067 n10__x1 vss 150.834e-18
c1068 n6__y1 vss 63.0729e-18
c1069 n18__x0 vss 287.985e-18
c1070 n14__y0 vss 197.628e-18
c1071 n24__vdd vss 3.62439e-18
c1072 n27__vdd vss 18.3439e-18
c1073 n28__vdd vss 39.4044e-18
c1074 n23__vdd vss 60.5487e-18
c1075 n39__clk4b vss 95.3292e-18
c1076 n15__y0 vss 226.792e-18
c1077 n14__y2 vss 477.552e-18
c1078 n17__x0 vss 242.443e-18
c1079 n14__x2 vss 353.096e-18
c1080 n66__clk4 vss 672.532e-18
c1081 n10__clkb vss 150.381e-18
c1082 n11__clkb vss 188.393e-18
c1083 n10__clk vss 14.5996e-18
c1084 n251__vddio vss 13.366e-18
c1085 n407__r_out vss 121.4e-18
c1086 n402__r_out vss 83.2188e-18
c1087 n249__vddio vss 105.951e-18
c1088 n396__r_out vss 100.572e-18
c1089 n398__r_out vss 128.828e-18
c1090 n245__vddio vss 100.945e-18
c1091 n388__r_out vss 101.019e-18
c1092 n390__r_out vss 128.974e-18
c1093 n241__vddio vss 101.019e-18
c1094 n380__r_out vss 100.823e-18
c1095 n382__r_out vss 128.779e-18
c1096 n237__vddio vss 100.462e-18
c1097 n372__r_out vss 100.462e-18
c1098 n374__r_out vss 128.641e-18
c1099 n233__vddio vss 100.823e-18
c1100 n364__r_out vss 101.019e-18
c1101 n366__r_out vss 128.974e-18
c1102 n229__vddio vss 101.019e-18
c1103 n356__r_out vss 100.823e-18
c1104 n358__r_out vss 128.779e-18
c1105 n225__vddio vss 100.462e-18
c1106 n348__r_out vss 100.462e-18
c1107 n350__r_out vss 128.641e-18
c1108 n221__vddio vss 100.823e-18
c1109 n340__r_out vss 101.019e-18
c1110 n342__r_out vss 128.974e-18
c1111 n217__vddio vss 101.019e-18
c1112 n332__r_out vss 100.823e-18
c1113 n334__r_out vss 128.779e-18
c1114 n213__vddio vss 100.462e-18
c1115 n324__r_out vss 100.462e-18
c1116 n326__r_out vss 128.641e-18
c1117 n209__vddio vss 100.282e-18
c1118 n316__r_out vss 100.282e-18
c1119 n318__r_out vss 128.204e-18
c1120 n205__vddio vss 96.3059e-18
c1121 n308__r_out vss 96.3059e-18
c1122 n310__r_out vss 125.682e-18
c1123 n201__vddio vss 96.537e-18
c1124 n300__r_out vss 96.44e-18
c1125 n302__r_out vss 127.033e-18
c1126 n197__vddio vss 97.3726e-18
c1127 n292__r_out vss 97.4712e-18
c1128 n294__r_out vss 127.953e-18
c1129 n193__vddio vss 96.8486e-18
c1130 n284__r_out vss 96.847e-18
c1131 n286__r_out vss 126.257e-18
c1132 n189__vddio vss 96.537e-18
c1133 n276__r_out vss 96.44e-18
c1134 n278__r_out vss 127.033e-18
c1135 n185__vddio vss 97.3726e-18
c1136 n268__r_out vss 97.4712e-18
c1137 n270__r_out vss 127.953e-18
c1138 n181__vddio vss 96.8486e-18
c1139 n260__r_out vss 96.847e-18
c1140 n262__r_out vss 126.257e-18
c1141 n177__vddio vss 96.537e-18
c1142 n252__r_out vss 96.44e-18
c1143 n254__r_out vss 127.033e-18
c1144 n173__vddio vss 97.3726e-18
c1145 n244__r_out vss 97.4712e-18
c1146 n246__r_out vss 127.953e-18
c1147 n169__vddio vss 96.8486e-18
c1148 n236__r_out vss 96.847e-18
c1149 n238__r_out vss 126.257e-18
c1150 n165__vddio vss 96.5018e-18
c1151 n228__r_out vss 96.4048e-18
c1152 n230__r_out vss 126.998e-18
c1153 n161__vddio vss 98.0275e-18
c1154 n220__r_out vss 98.3219e-18
c1155 n222__r_out vss 128.838e-18
c1156 n157__vddio vss 101.608e-18
c1157 n212__r_out vss 101.411e-18
c1158 n214__r_out vss 129.658e-18
c1159 n153__vddio vss 100.898e-18
c1160 n204__r_out vss 101.094e-18
c1161 n206__r_out vss 129.049e-18
c1162 n149__vddio vss 97.0744e-18
c1163 n196__r_out vss 96.8787e-18
c1164 n198__r_out vss 126.291e-18
c1165 n145__vddio vss 100.38e-18
c1166 n188__r_out vss 100.024e-18
c1167 n190__r_out vss 128.558e-18
c1168 n141__vddio vss 100.768e-18
c1169 n184__r_out vss 97.2002e-18
c1170 n178__r_out vss 129.049e-18
c1171 n136__vddio vss 161.036e-18
c1172 n172__r_out vss 97.3625e-18
c1173 n174__r_out vss 126.291e-18
c1174 n132__vddio vss 100.38e-18
c1175 n164__r_out vss 100.38e-18
c1176 n166__r_out vss 128.558e-18
c1177 n128__vddio vss 100.898e-18
c1178 n156__r_out vss 101.094e-18
c1179 n158__r_out vss 129.049e-18
c1180 n124__vddio vss 97.0744e-18
c1181 n148__r_out vss 96.8787e-18
c1182 n150__r_out vss 126.291e-18
c1183 n120__vddio vss 100.38e-18
c1184 n140__r_out vss 100.38e-18
c1185 n142__r_out vss 128.558e-18
c1186 n116__vddio vss 100.357e-18
c1187 n132__r_out vss 100.357e-18
c1188 n134__r_out vss 128.279e-18
c1189 n112__vddio vss 100.266e-18
c1190 n124__r_out vss 100.266e-18
c1191 n126__r_out vss 128.188e-18
c1192 n108__vddio vss 96.4266e-18
c1193 n116__r_out vss 96.4266e-18
c1194 n118__r_out vss 126.063e-18
c1195 n104__vddio vss 97.4119e-18
c1196 n108__r_out vss 97.5106e-18
c1197 n110__r_out vss 127.885e-18
c1198 n100__vddio vss 100.906e-18
c1199 n100__r_out vss 100.807e-18
c1200 n102__r_out vss 128.763e-18
c1201 n96__vddio vss 96.4266e-18
c1202 n92__r_out vss 96.4266e-18
c1203 n94__r_out vss 126.063e-18
c1204 n92__vddio vss 97.8407e-18
c1205 n84__r_out vss 98.0699e-18
c1206 n86__r_out vss 128.467e-18
c1207 n88__vddio vss 101.483e-18
c1208 n76__r_out vss 101.254e-18
c1209 n78__r_out vss 129.232e-18
c1210 n84__vddio vss 100.462e-18
c1211 n68__r_out vss 100.462e-18
c1212 n70__r_out vss 128.641e-18
c1213 n80__vddio vss 100.823e-18
c1214 n60__r_out vss 101.019e-18
c1215 n62__r_out vss 128.974e-18
c1216 n76__vddio vss 101.019e-18
c1217 n52__r_out vss 100.823e-18
c1218 n54__r_out vss 128.779e-18
c1219 n72__vddio vss 100.462e-18
c1220 n44__r_out vss 100.462e-18
c1221 n46__r_out vss 128.641e-18
c1222 n68__vddio vss 100.643e-18
c1223 n36__r_out vss 100.773e-18
c1224 n38__r_out vss 128.718e-18
c1225 n64__vddio vss 100.813e-18
c1226 n28__r_out vss 100.878e-18
c1227 n30__r_out vss 128.856e-18
c1228 n60__vddio vss 97.0744e-18
c1229 n20__r_out vss 96.8787e-18
c1230 n22__r_out vss 126.291e-18
c1231 n56__vddio vss 99.456e-18
c1232 n12__r_out vss 100.379e-18
c1233 n14__r_out vss 128.597e-18
c1234 n52__vddio vss 246.362e-18
c1235 n4__r_out vss 72.9667e-18
c1236 n6__r_out vss 102.829e-18
c1237 n90__i12__net3 vss 79.0625e-18
c1238 n95__i12__net3 vss 93.8489e-18
c1239 n45__vddio vss 94.5797e-18
c1240 n78__i12__net3 vss 166.63e-18
c1241 n81__i12__net3 vss 141.349e-18
c1242 n41__vddio vss 105.555e-18
c1243 n62__i12__net3 vss 166.359e-18
c1244 n65__i12__net3 vss 142.031e-18
c1245 n37__vddio vss 106.515e-18
c1246 n46__i12__net3 vss 167.028e-18
c1247 n49__i12__net3 vss 141.336e-18
c1248 n33__vddio vss 105.699e-18
c1249 n30__i12__net3 vss 165.929e-18
c1250 n33__i12__net3 vss 141.395e-18
c1251 n29__vddio vss 105.647e-18
c1252 n14__i12__net3 vss 157.51e-18
c1253 n17__i12__net3 vss 131.314e-18
c1254 n19__vddio vss 75.1303e-18
c1255 n41__i12__net2 vss 80.8265e-18
c1256 n42__i12__net2 vss 80.4634e-18
c1257 n24__vddio vss 115.847e-18
c1258 n34__i12__net2 vss 111.71e-18
c1259 n37__i12__net2 vss 74.3787e-18
c1260 n270__vdd vss 24.7385e-18
c1261 n7__i11__net1 vss 25.0687e-18
c1262 n5__i11__net1 vss 58.1358e-18
c1263 n6__vddio vss 8.00573e-18
c1264 n9__i14__i5__net5 vss 64.3599e-18
c1265 n39__clk vss 211.409e-18
c1266 n13__r0 vss 49.6945e-18
c1267 n37__i14__shift vss 130.561e-18
c1268 n26__clkb vss 224.553e-18
c1269 n8__i14__net14 vss 79.0844e-18
c1270 n5__i14__net14 vss 92.3745e-18
c1271 n5__i14__i5__net5 vss 176.728e-18
c1272 n36__i14__shift vss 166.494e-18
c1273 n5__i14__i2__net1 vss 94.7583e-18
c1274 n38__clk vss 180.997e-18
c1275 n8__i14__net15 vss 76.89e-18
c1276 n7__serial_out vss 124.42e-18
c1277 n6__i14__i2__net1 vss 147.37e-18
c1278 n35__i14__shift vss 124.057e-18
c1279 n9__r1 vss 156.439e-18
c1280 n70__rst vss 98.5499e-18
c1281 n265__vdd vss 81.1369e-18
c1282 n34__i14__shift vss 121.858e-18
c1283 n6__i14__net8 vss 97.5755e-18
c1284 n9__i14__i4__net5 vss 115.112e-18
c1285 n33__i14__shift vss 163.809e-18
c1286 n5__i14__i1__net1 vss 119.597e-18
c1287 n4__i14__net8 vss 89.0317e-18
c1288 n8__i14__net9 vss 76.6252e-18
c1289 n36__clk vss 246.629e-18
c1290 n8__i14__i1__net1 vss 145.431e-18
c1291 n25__clkb vss 141.798e-18
c1292 n251__vdd vss 243.625e-18
c1293 n32__i14__shift vss 129.124e-18
c1294 n5__i14__i4__net5 vss 204.22e-18
c1295 n35__clk vss 160.968e-18
c1296 n7__r2 vss 131.691e-18
c1297 n31__i14__shift vss 130.026e-18
c1298 n2__i14__net15 vss 133.167e-18
c1299 n6__i14__net2 vss 87.0354e-18
c1300 n7__i14__net2 vss 114.432e-18
c1301 n30__i14__shift vss 141.01e-18
c1302 n5__i14__i0__net1 vss 122.452e-18
c1303 n248__vdd vss 86.1883e-18
c1304 n6__i14__i0__net1 vss 126.112e-18
c1305 n29__i14__shift vss 124.484e-18
c1306 n9__i14__i3__net5 vss 119.229e-18
c1307 n29__clk vss 146.367e-18
c1308 n24__clkb vss 140.876e-18
c1309 n232__vdd vss 143.156e-18
c1310 n5__i14__i3__net5 vss 203.322e-18
c1311 n234__vdd vss 74.8323e-18
c1312 n236__vdd vss 21.7181e-18
c1313 n231__vdd vss 113.346e-18
c1314 n27__clk vss 170.145e-18
c1315 n2__i14__net9 vss 184.544e-18
c1316 n25__i14__shift vss 83.2204e-18
c1317 n9__i14__i7__net1 vss 83.3681e-18
c1318 n63__rst vss 88.758e-18
c1319 n8__i14__i7__net1 vss 77.6556e-18
c1320 n20__clk2 vss 489.392e-18
c1321 n6__i14__i7__net1 vss 104.059e-18
c1322 n72__clk4 vss 387.518e-18
c1323 n4__r1 vss 60.1965e-18
c1324 n5__r1 vss 60.471e-18
c1325 n19__i10__net116 vss 202.301e-18
c1326 n2__r1 vss 102.046e-18
c1327 n16__i10__net114 vss 86.2244e-18
c1328 n17__i10__net114 vss 93.3308e-18
c1329 n14__i10__net114 vss 126.639e-18
c1330 n12__i10__net114 vss 55.1366e-18
c1331 n18__s1 vss 155.122e-18
c1332 n186__vdd vss 23.4559e-18
c1333 n187__vdd vss 24.825e-18
c1334 n4__i10__net125 vss 113.141e-18
c1335 n17__s0 vss 217.153e-18
c1336 n4__i10__net122 vss 47.7198e-18
c1337 n15__net12 vss 205.076e-18
c1338 n9__i10__net114 vss 111.874e-18
c1339 n8__i10__net114 vss 92.5684e-18
c1340 n18__i10__net116 vss 275.367e-18
c1341 n2__r0 vss 166.736e-18
c1342 n9__i9__net51 vss 143.336e-18
c1343 n2__i10__net115 vss 106.564e-18
c1344 n2__i10__net124 vss 55.1256e-18
c1345 n16__s1 vss 54.4241e-18
c1346 n4__i9__net51 vss 135.062e-18
c1347 n9__i10__net116 vss 43.5232e-18
c1348 n10__i10__net116 vss 160.086e-18
c1349 n14__s0 vss 304.352e-18
c1350 n20__c1 vss 191.026e-18
c1351 n17__net12 vss 419.349e-18
c1352 n21__c0 vss 215.936e-18
c1353 n15__a1 vss 223.931e-18
c1354 n14__a3 vss 164.073e-18
c1355 n16__a0 vss 217.895e-18
c1356 n16__a2 vss 220.304e-18
c1357 n19__c0 vss 104.374e-18
c1358 n18__c1 vss 165.074e-18
c1359 n10__s0 vss 278.001e-18
c1360 n10__s1 vss 160.374e-18
c1361 n9__i7__net51 vss 113.234e-18
c1362 n9__i8__net51 vss 94.0622e-18
c1363 n151__vdd vss 25.4868e-18
c1364 n148__vdd vss 44.6468e-18
c1365 n13__a1 vss 428.158e-18
c1366 n13__a3 vss 308.243e-18
c1367 n4__i7__net51 vss 122.91e-18
c1368 n4__i8__net51 vss 122.675e-18
c1369 n13__a0 vss 591.011e-18
c1370 n13__a2 vss 578.295e-18
c1371 n9__a3 vss 219.979e-18
c1372 n12__a1 vss 175.165e-18
c1373 n23__y1 vss 60.7267e-18
c1374 n15__i1__rstb vss 225.578e-18
c1375 n15__i2__rstb vss 233.769e-18
c1376 n43__rst vss 95.6363e-18
c1377 n36__rst vss 104.971e-18
c1378 n11__i1__net4 vss 261.694e-18
c1379 n11__i2__net4 vss 275.398e-18
c1380 n14__y3 vss 86.5049e-18
c1381 n22__x1 vss 51.1378e-18
c1382 n60__clk4 vss 140.503e-18
c1383 n59__clk4 vss 139.368e-18
c1384 n79__vdd vss 186.761e-18
c1385 n73__vdd vss 67.7587e-18
c1386 n8__i1__net2 vss 171.429e-18
c1387 n8__i2__net2 vss 179.612e-18
c1388 n11__y3 vss 115.18e-18
c1389 n46__clk4b vss 258.546e-18
c1390 n45__clk4b vss 246.51e-18
c1391 n20__y1 vss 80.9585e-18
c1392 n78__vdd vss 124.729e-18
c1393 n71__vdd vss 62.5195e-18
c1394 n58__clk4 vss 339.415e-18
c1395 n68__vdd vss 21.3697e-18
c1396 n57__clk4 vss 332.669e-18
c1397 n66__vdd vss 76.7531e-18
c1398 n19__x1 vss 88.7945e-18
c1399 n11__x3 vss 53.2184e-18
c1400 n6__i1__net2 vss 141.317e-18
c1401 n6__i2__net2 vss 139.352e-18
c1402 n65__vdd vss 164.893e-18
c1403 n64__vdd vss 67.6557e-18
c1404 n11__i1__rstb vss 35.7041e-18
c1405 n11__i2__rstb vss 107.108e-18
c1406 n9__y3 vss 189.586e-18
c1407 n30__rst vss 83.9473e-18
c1408 n29__rst vss 107.115e-18
c1409 n16__x2 vss 180.073e-18
c1410 n16__y2 vss 178.586e-18
c1411 n62__vdd vss 61.8975e-18
c1412 n8__x3 vss 135.675e-18
c1413 n54__clk4 vss 192.955e-18
c1414 n51__clk4 vss 191.643e-18
c1415 n9__i1__net4 vss 288.434e-18
c1416 n9__i2__net4 vss 233.436e-18
c1417 n44__clk4b vss 127.938e-18
c1418 n43__clk4b vss 126.838e-18
c1419 n50__clk4 vss 238.816e-18
c1420 n49__clk4 vss 241.185e-18
c1421 n6__i1__net4 vss 97.0185e-18
c1422 n6__i2__net4 vss 109.1e-18
c1423 n11__x1 vss 82.3778e-18
c1424 n11__y1 vss 83.4796e-18
c1425 n48__clk4 vss 148.993e-18
c1426 n47__clk4 vss 149.373e-18
c1427 n8__i1__net3 vss 144.945e-18
c1428 n8__i2__net3 vss 152.003e-18
c1429 n42__clk4b vss 121.719e-18
c1430 n41__clk4b vss 121.831e-18
c1431 n46__clk4 vss 298.973e-18
c1432 n45__clk4 vss 313.77e-18
c1433 n4__a0 vss 288.288e-18
c1434 n6__i1__net3 vss 107.567e-18
c1435 n6__i2__net3 vss 112.065e-18
c1436 n4__a2 vss 438.754e-18
c1437 n9__i1__rstb vss 309.054e-18
c1438 n9__i2__rstb vss 306.445e-18
c1439 n17__y0 vss 113.599e-18
c1440 n10__i1__net1 vss 88.1008e-18
c1441 n10__i2__net1 vss 90.3447e-18
c1442 n20__rst vss 107.619e-18
c1443 n19__rst vss 107.165e-18
c1444 n11__y2 vss 61.198e-18
c1445 n9__x1 vss 51.6346e-18
c1446 n5__y1 vss 142.108e-18
c1447 n18__rst vss 129.476e-18
c1448 n17__rst vss 123.705e-18
c1449 n10__y0 vss 67.2241e-18
c1450 n11__x0 vss 54.1966e-18
c1451 n31__vdd vss 163.72e-18
c1452 n21__vdd vss 78.0673e-18
c1453 n44__clk4 vss 137.323e-18
c1454 n43__clk4 vss 140.721e-18
c1455 n8__i1__net1 vss 175.148e-18
c1456 n8__i2__net1 vss 185.348e-18
c1457 n11__x2 vss 52.6933e-18
c1458 n30__vdd vss 162.659e-18
c1459 n19__vdd vss 65.2347e-18
c1460 n25__vdd vss 48.5503e-18
c1461 n26__vdd vss 24.5112e-18
c1462 n29__vdd vss 150.496e-18
c1463 n22__vdd vss 170.29e-18
c1464 n38__clk4b vss 301.017e-18
c1465 n37__clk4b vss 269.056e-18
c1466 n9__y0 vss 80.9817e-18
c1467 n17__vdd vss 68.1404e-18
c1468 n9__y2 vss 80.9754e-18
c1469 n42__clk4 vss 203.889e-18
c1470 n41__clk4 vss 222.381e-18
c1471 n8__x0 vss 138.258e-18
c1472 n15__vdd vss 62.8902e-18
c1473 n8__x2 vss 86.934e-18
c1474 n6__i1__net1 vss 86.6049e-18
c1475 n6__i2__net1 vss 84.4899e-18
c1476 n32__clk4b vss 215.96e-18
c1477 n34__clk4 vss 175.155e-18
c1478 n11__i0__net4 vss 103.219e-18
c1479 n15__clk2 vss 141.635e-18
c1480 n9__i0__net6 vss 122.119e-18
c1481 n9__i0__net4 vss 125.218e-18
c1482 n16__i0__net1 vss 177.192e-18
c1483 n14__clk2 vss 164.184e-18
c1484 n6__i0__net6 vss 108.751e-18
c1485 n13__clk2 vss 819.656e-18
c1486 n13__i0__net1 vss 129.37e-18
c1487 n11__i0__net1 vss 133.603e-18
c1488 n10__clk2 vss 89.1792e-18
c1489 n6__clkb vss 10.4505e-18
c1490 n13__clk vss 153.966e-18
c1491 n9__i0__net2 vss 137.18e-18
c1492 n9__i0__net1 vss 119.379e-18
c1493 n11__clk vss 295.02e-18
c1494 n1__vdd vss 7.8169e-18
c1495 n6__i0__net2 vss 87.258e-18
c1496 n12__clk vss 152.694e-18
c1497 n13__vddio vss 28.4106e-15
c1498 n403__r_out vss 357.414e-18
c1499 n399__r_out vss 428.183e-18
c1500 n391__r_out vss 426.363e-18
c1501 n383__r_out vss 426.913e-18
c1502 n375__r_out vss 426.645e-18
c1503 n367__r_out vss 426.363e-18
c1504 n359__r_out vss 426.913e-18
c1505 n351__r_out vss 426.645e-18
c1506 n343__r_out vss 426.363e-18
c1507 n335__r_out vss 426.913e-18
c1508 n327__r_out vss 426.645e-18
c1509 n319__r_out vss 426.82e-18
c1510 n311__r_out vss 427.954e-18
c1511 n303__r_out vss 427.886e-18
c1512 n295__r_out vss 427.805e-18
c1513 n287__r_out vss 427.954e-18
c1514 n279__r_out vss 427.886e-18
c1515 n271__r_out vss 427.805e-18
c1516 n263__r_out vss 427.954e-18
c1517 n255__r_out vss 427.886e-18
c1518 n247__r_out vss 427.805e-18
c1519 n239__r_out vss 427.954e-18
c1520 n231__r_out vss 427.961e-18
c1521 n223__r_out vss 427.321e-18
c1522 n215__r_out vss 426.633e-18
c1523 n207__r_out vss 426.14e-18
c1524 n199__r_out vss 428.262e-18
c1525 n191__r_out vss 426.644e-18
c1526 n179__r_out vss 426.159e-18
c1527 n405__r_out vss 686.708e-18
c1528 n247__vddio vss 974.949e-18
c1529 n393__r_out vss 967.711e-18
c1530 n243__vddio vss 958.246e-18
c1531 n385__r_out vss 963.93e-18
c1532 n239__vddio vss 957.696e-18
c1533 n377__r_out vss 964.48e-18
c1534 n235__vddio vss 958.246e-18
c1535 n369__r_out vss 964.48e-18
c1536 n231__vddio vss 958.246e-18
c1537 n361__r_out vss 963.93e-18
c1538 n227__vddio vss 957.696e-18
c1539 n353__r_out vss 964.48e-18
c1540 n223__vddio vss 958.246e-18
c1541 n345__r_out vss 964.48e-18
c1542 n219__vddio vss 958.246e-18
c1543 n337__r_out vss 963.93e-18
c1544 n215__vddio vss 957.696e-18
c1545 n329__r_out vss 964.48e-18
c1546 n211__vddio vss 958.246e-18
c1547 n321__r_out vss 964.48e-18
c1548 n207__vddio vss 958.246e-18
c1549 n313__r_out vss 964.387e-18
c1550 n203__vddio vss 960.835e-18
c1551 n305__r_out vss 966.862e-18
c1552 n199__vddio vss 960.532e-18
c1553 n297__r_out vss 967.062e-18
c1554 n195__vddio vss 960.731e-18
c1555 n289__r_out vss 966.713e-18
c1556 n191__vddio vss 960.673e-18
c1557 n281__r_out vss 966.862e-18
c1558 n187__vddio vss 960.532e-18
c1559 n273__r_out vss 967.062e-18
c1560 n183__vddio vss 960.731e-18
c1561 n265__r_out vss 966.713e-18
c1562 n179__vddio vss 960.673e-18
c1563 n257__r_out vss 966.862e-18
c1564 n175__vddio vss 960.532e-18
c1565 n249__r_out vss 967.062e-18
c1566 n171__vddio vss 960.731e-18
c1567 n241__r_out vss 966.713e-18
c1568 n167__vddio vss 960.673e-18
c1569 n233__r_out vss 966.862e-18
c1570 n163__vddio vss 960.532e-18
c1571 n225__r_out vss 967.137e-18
c1572 n159__vddio vss 960.806e-18
c1573 n217__r_out vss 966.229e-18
c1574 n155__vddio vss 957.507e-18
c1575 n209__r_out vss 964.468e-18
c1576 n151__vddio vss 958.234e-18
c1577 n201__r_out vss 963.707e-18
c1578 n147__vddio vss 960.155e-18
c1579 n193__r_out vss 967.17e-18
c1580 n143__vddio vss 958.258e-18
c1581 n185__r_out vss 964.479e-18
c1582 n139__vddio vss 958.633e-18
c1583 n181__r_out vss 966.327e-18
c1584 n134__vddio vss 853.255e-18
c1585 n169__r_out vss 969.183e-18
c1586 n130__vddio vss 958.324e-18
c1587 n161__r_out vss 964.479e-18
c1588 n126__vddio vss 958.246e-18
c1589 n153__r_out vss 963.707e-18
c1590 n122__vddio vss 960.155e-18
c1591 n145__r_out vss 967.17e-18
c1592 n118__vddio vss 958.255e-18
c1593 n137__r_out vss 964.479e-18
c1594 n114__vddio vss 958.246e-18
c1595 n129__r_out vss 964.379e-18
c1596 n110__vddio vss 958.145e-18
c1597 n121__r_out vss 964.487e-18
c1598 n106__vddio vss 960.935e-18
c1599 n113__r_out vss 966.865e-18
c1600 n102__vddio vss 960.534e-18
c1601 n105__r_out vss 966.713e-18
c1602 n98__vddio vss 957.894e-18
c1603 n97__r_out vss 964.487e-18
c1604 n94__vddio vss 960.935e-18
c1605 n89__r_out vss 966.934e-18
c1606 n90__vddio vss 960.603e-18
c1607 n81__r_out vss 966.411e-18
c1608 n86__vddio vss 957.592e-18
c1609 n73__r_out vss 964.55e-18
c1610 n82__vddio vss 958.316e-18
c1611 n65__r_out vss 964.48e-18
c1612 n78__vddio vss 958.246e-18
c1613 n57__r_out vss 963.93e-18
c1614 n74__vddio vss 957.696e-18
c1615 n49__r_out vss 964.48e-18
c1616 n70__vddio vss 958.246e-18
c1617 n41__r_out vss 964.48e-18
c1618 n66__vddio vss 958.246e-18
c1619 n33__r_out vss 964.019e-18
c1620 n62__vddio vss 957.785e-18
c1621 n25__r_out vss 963.649e-18
c1622 n58__vddio vss 960.097e-18
c1623 n17__r_out vss 968.666e-18
c1624 n54__vddio vss 958.253e-18
c1625 n9__r_out vss 975.622e-18
c1626 n50__vddio vss 933.357e-18
c1627 n1__r_out vss 810.389e-18
c1628 n361__i12__net3 vss 731.25e-18
c1629 n42__vddio vss 982.722e-18
c1630 n74__i12__net3 vss 920.134e-18
c1631 n38__vddio vss 966.913e-18
c1632 n58__i12__net3 vss 918.488e-18
c1633 n34__vddio vss 967.101e-18
c1634 n42__i12__net3 vss 918.205e-18
c1635 n30__vddio vss 967.266e-18
c1636 n26__i12__net3 vss 918.87e-18
c1637 n26__vddio vss 968.636e-18
c1638 n10__i12__net3 vss 927.404e-18
c1639 n15__vddio vss 631.614e-18
c1640 n43__i12__net2 vss 430.187e-18
c1641 n21__vddio vss 761.912e-18
c1642 n31__i12__net2 vss 407.33e-18
c1643 n7__i12__net1 vss 147.947e-18
c1644 n175__r_out vss 430.323e-18
c1645 n167__r_out vss 426.644e-18
c1646 n159__r_out vss 426.14e-18
c1647 n151__r_out vss 428.262e-18
c1648 n143__r_out vss 426.644e-18
c1649 n135__r_out vss 426.812e-18
c1650 n127__r_out vss 426.92e-18
c1651 n119__r_out vss 427.689e-18
c1652 n111__r_out vss 427.805e-18
c1653 n103__r_out vss 426.92e-18
c1654 n95__r_out vss 427.758e-18
c1655 n87__r_out vss 427.503e-18
c1656 n79__r_out vss 426.983e-18
c1657 n71__r_out vss 426.645e-18
c1658 n63__r_out vss 426.363e-18
c1659 n55__r_out vss 426.913e-18
c1660 n47__r_out vss 426.645e-18
c1661 n39__r_out vss 426.452e-18
c1662 n31__r_out vss 426.082e-18
c1663 n23__r_out vss 429.157e-18
c1664 n15__r_out vss 432.757e-18
c1665 n7__r_out vss 358.931e-18
c1666 n366__i12__net3 vss 374.681e-18
c1667 n82__i12__net3 vss 432.837e-18
c1668 n66__i12__net3 vss 431.424e-18
c1669 n50__i12__net3 vss 432.237e-18
c1670 n34__i12__net3 vss 431.807e-18
c1671 n18__i12__net3 vss 437.733e-18
c1672 n47__i12__net2 vss 208.267e-18
c1673 n36__i12__net2 vss 193.655e-18
c1674 n9__i12__net1 vss 87.1732e-18
c1675 n272__vdd vss 47.5304e-18
c1676 n4__vddio vss 166.693e-18
c1677 n25__vddio vss 242.349e-18
c1678 n9__r_in vss 178.682e-18
c1679 n6__i11__net1 vss 53.9803e-18
c1680 n4__net5 vss 236.956e-18
c1681 n274__vdd vss 39.0235e-18
c1682 n6__r_in vss 74.1696e-18
c1683 n2__vddio vss 62.7164e-18
c1684 n5__net5 vss 75.6929e-18
c1685 n6__i14__i5__net5 vss 69.6988e-18
c1686 n11__r0 vss 90.498e-18
c1687 n268__vdd vss 182.221e-18
c1688 n4__i14__net14 vss 52.0767e-18
c1689 n7__i14__net15 vss 64.8173e-18
c1690 n6__serial_out vss 64.5135e-18
c1691 n9__i14__i2__net1 vss 48.2126e-18
c1692 n4__i14__i5__net5 vss 96.3678e-18
c1693 n253__vdd vss 83.8994e-18
c1694 n8__i14__i5__net5 vss 77.9854e-18
c1695 n10__r0 vss 73.3781e-18
c1696 n6__i14__net14 vss 77.6908e-18
c1697 n9__i14__net15 vss 76.9325e-18
c1698 n8__serial_out vss 36.3051e-18
c1699 n7__i14__i2__net1 vss 81.841e-18
c1700 n10__serial_out vss 38.6525e-18
c1701 n254__vdd vss 384.404e-18
c1702 n229__vdd vss 545.525e-18
c1703 n10__r1 vss 103.283e-18
c1704 n4__i14__i5__rstb vss 57.3162e-18
c1705 n266__vdd vss 71.1675e-18
c1706 n8__r1 vss 48.0007e-18
c1707 n5__i14__i5__rstb vss 51.8668e-18
c1708 n5__i14__net8 vss 52.4878e-18
c1709 n6__i14__i4__net5 vss 79.2265e-18
c1710 n7__i14__net9 vss 66.2158e-18
c1711 n9__i14__i1__net1 vss 53.8052e-18
c1712 n252__vdd vss 68.6993e-18
c1713 n258__vdd vss 75.1426e-18
c1714 n6__r2 vss 47.2622e-18
c1715 n8__i14__net2 vss 52.8545e-18
c1716 n4__i14__i4__net5 vss 98.6607e-18
c1717 n7__i14__net8 vss 78.3785e-18
c1718 n8__i14__i4__net5 vss 90.4437e-18
c1719 n9__i14__net9 vss 77.6173e-18
c1720 n6__i14__i1__net1 vss 90.755e-18
c1721 n8__r2 vss 103.64e-18
c1722 n3__i14__net15 vss 41.6096e-18
c1723 n9__i14__net2 vss 76.8005e-18
c1724 n5__i14__net15 vss 38.9934e-18
c1725 n7__i14__i0__net1 vss 84.6623e-18
c1726 n4__i14__i4__rstb vss 59.4079e-18
c1727 n249__vdd vss 72.1501e-18
c1728 n9__i14__i0__net1 vss 50.7972e-18
c1729 n5__i14__i4__rstb vss 53.8012e-18
c1730 n259__vdd vss 49.5621e-18
c1731 n6__i14__i3__net5 vss 78.9509e-18
c1732 n233__vdd vss 69.0506e-18
c1733 n28__i14__shift vss 41.2809e-18
c1734 n4__i14__i3__net5 vss 96.1305e-18
c1735 n8__i14__i3__net5 vss 90.2156e-18
c1736 n3__i14__net9 vss 41.0046e-18
c1737 n261__vdd vss 119.262e-18
c1738 n27__i14__shift vss 35.0658e-18
c1739 n5__i14__net9 vss 38.923e-18
c1740 n263__vdd vss 62.6775e-18
c1741 n228__vdd vss 71.7989e-18
c1742 n7__i14__i7__net1 vss 61.741e-18
c1743 n5__i14__i3__rstb vss 42.9708e-18
c1744 n264__vdd vss 89.1172e-18
c1745 n4__i14__i3__rstb vss 51.9585e-18
c1746 n165__vdd vss 819.634e-18
c1747 n4__r2 vss 80.2253e-18
c1748 n217__vdd vss 70.6869e-18
c1749 n218__vdd vss 64.1798e-18
c1750 n219__vdd vss 78.6188e-18
c1751 n11__i10__net114 vss 79.1509e-18
c1752 n191__vdd vss 37.7906e-18
c1753 n220__vdd vss 107.297e-18
c1754 n4__i9__carry_bar vss 103.46e-18
c1755 n7__i10__net122 vss 166.593e-21
c1756 n200__vdd vss 40.1266e-18
c1757 n221__vdd vss 127.131e-18
c1758 n201__vdd vss 40.525e-18
c1759 n2__i10__net122 vss 58.0245e-18
c1760 n13__net12 vss 137.748e-18
c1761 n7__i10__net114 vss 107.227e-18
c1762 n7__i10__net115 vss 94.7375e-18
c1763 n222__vdd vss 192.769e-18
c1764 n3__i10__net115 vss 99.6318e-18
c1765 n202__vdd vss 97.5332e-18
c1766 n8__i9__net51 vss 46.2761e-18
c1767 n11__i10__net116 vss 126.346e-18
c1768 n2__i9__net49 vss 166.018e-18
c1769 n203__vdd vss 56.7794e-18
c1770 n198__vdd vss 52.4068e-18
c1771 n13__i10__net116 vss 62.2145e-18
c1772 n223__vdd vss 97.7179e-18
c1773 n3__r2 vss 34.7071e-18
c1774 n3__r1 vss 56.9673e-18
c1775 n13__i10__net114 vss 60.1342e-18
c1776 n5__i10__net125 vss 68.553e-21
c1777 n6__i9__carry_bar vss 102.933e-18
c1778 n16__net12 vss 132.027e-18
c1779 n10__i10__net114 vss 76.937e-18
c1780 n8__i10__net124 vss 54.258e-18
c1781 n5__r0 vss 35.344e-18
c1782 n3__i10__net124 vss 63.5774e-18
c1783 n14__i10__net116 vss 79.6249e-18
c1784 n4__r0 vss 95.0503e-18
c1785 n17__i10__net116 vss 41.5213e-18
c1786 n180__vdd vss 965.624e-18
c1787 n167__vdd vss 67.4189e-18
c1788 n152__vdd vss 51.901e-18
c1789 n4__i7__carry_bar vss 108.461e-18
c1790 n4__i8__carry_bar vss 105.994e-18
c1791 n176__vdd vss 41.5641e-18
c1792 n161__vdd vss 40.7557e-18
c1793 n177__vdd vss 42.1432e-18
c1794 n162__vdd vss 36.5755e-18
c1795 n17__c0 vss 140.635e-18
c1796 n17__c1 vss 141.961e-18
c1797 n9__s0 vss 120.032e-18
c1798 n9__s1 vss 121.261e-18
c1799 n178__vdd vss 99.1438e-18
c1800 n8__i7__net51 vss 45.2817e-18
c1801 n163__vdd vss 93.8445e-18
c1802 n8__i8__net51 vss 45.5453e-18
c1803 n2__i7__net49 vss 166.081e-18
c1804 n2__i8__net49 vss 166.223e-18
c1805 n179__vdd vss 56.087e-18
c1806 n174__vdd vss 53.0187e-18
c1807 n164__vdd vss 55.0681e-18
c1808 n159__vdd vss 51.038e-18
c1809 n6__i7__carry_bar vss 104.47e-18
c1810 n6__i8__carry_bar vss 106.298e-18
c1811 n20__c0 vss 132.692e-18
c1812 n19__c1 vss 40.6008e-18
c1813 n13__s0 vss 35.2155e-18
c1814 n13__s1 vss 35.8761e-18
c1815 n12__s0 vss 99.0057e-18
c1816 n12__s1 vss 97.6862e-18
c1817 n138__vdd vss 138.555e-18
c1818 n13__i1__rstb vss 42.1929e-18
c1819 n13__i2__rstb vss 38.6439e-18
c1820 n111__vdd vss 118.317e-18
c1821 n96__vdd vss 125.419e-18
c1822 n9__a1 vss 106.225e-18
c1823 n13__i1__net4 vss 58.2089e-18
c1824 n13__i2__net4 vss 57.8557e-18
c1825 n19__x3 vss 83.7949e-18
c1826 n19__y3 vss 83.3123e-18
c1827 n74__vdd vss 118.123e-18
c1828 n72__vdd vss 67.1881e-18
c1829 n119__vdd vss 92.0928e-18
c1830 n104__vdd vss 90.2996e-18
c1831 n4__i4__bbar vss 163.056e-18
c1832 n12__a3 vss 103.134e-18
c1833 n70__vdd vss 59.515e-18
c1834 n4__i4__abar vss 243.059e-18
c1835 n4__i1__net2 vss 99.1897e-18
c1836 n4__i2__net2 vss 99.8135e-18
c1837 n63__vdd vss 66.6273e-18
c1838 n120__vdd vss 77.3097e-18
c1839 n105__vdd vss 77.5363e-18
c1840 n4__i6__bbar vss 167.145e-18
c1841 n16__i1__rstb vss 45.0997e-18
c1842 n16__i2__rstb vss 45.582e-18
c1843 n16__x3 vss 47.5783e-18
c1844 n16__y3 vss 47.8086e-18
c1845 n11__a1 vss 92.7839e-18
c1846 n17__x3 vss 88.8605e-18
c1847 n17__y3 vss 88.5846e-18
c1848 n2__i4__net3 vss 131.004e-18
c1849 n6__i4__bbar vss 124.083e-18
c1850 n11__a3 vss 95.5817e-18
c1851 n6__i4__abar vss 117.035e-18
c1852 n7__i1__net2 vss 82.2372e-18
c1853 n7__i2__net2 vss 84.4876e-18
c1854 n2__i6__net3 vss 134.104e-18
c1855 n139__vdd vss 152.895e-18
c1856 n6__i6__bbar vss 126.037e-18
c1857 n124__vdd vss 786.015e-18
c1858 n109__vdd vss 355.675e-18
c1859 n76__vdd vss 176.505e-18
c1860 n15__x2 vss 62.6992e-18
c1861 n15__y2 vss 64.4638e-18
c1862 n6__i6__abar vss 114.689e-18
c1863 n17__x2 vss 47.7725e-18
c1864 n17__y2 vss 48.8721e-18
c1865 n61__vdd vss 60.0479e-18
c1866 n4__i6__abar vss 248.433e-18
c1867 n121__vdd vss 91.9802e-18
c1868 n106__vdd vss 91.9937e-18
c1869 n7__i1__net4 vss 104.993e-18
c1870 n7__i2__net4 vss 104.809e-18
c1871 n16__x1 vss 27.2603e-18
c1872 n16__y1 vss 27.6611e-18
c1873 n7__i1__net3 vss 88.2903e-18
c1874 n7__i2__net3 vss 88.4791e-18
c1875 n8__x1 vss 42.4073e-18
c1876 n4__y1 vss 44.417e-18
c1877 n60__vdd vss 174.945e-18
c1878 n57__vdd vss 154.559e-18
c1879 n4__i1__net4 vss 82.1325e-18
c1880 n4__i2__net4 vss 81.4472e-18
c1881 n15__x1 vss 64.3919e-18
c1882 n15__y1 vss 63.889e-18
c1883 n122__vdd vss 89.4676e-18
c1884 n107__vdd vss 89.5252e-18
c1885 n4__i1__net3 vss 100.816e-18
c1886 n4__i2__net3 vss 101.198e-18
c1887 n123__vdd vss 92.7527e-18
c1888 n108__vdd vss 92.5633e-18
c1889 n58__vdd vss 129.205e-18
c1890 n55__vdd vss 115.757e-18
c1891 n9__i1__net1 vss 61.6458e-18
c1892 n9__i2__net1 vss 61.6678e-18
c1893 n14__x0 vss 85.1874e-18
c1894 n11__y0 vss 85.6579e-18
c1895 n20__vdd vss 70.28e-18
c1896 n18__vdd vss 74.1916e-18
c1897 n4__i3__bbar vss 161.957e-18
c1898 n125__vdd vss 79.1e-18
c1899 n110__vdd vss 79.5244e-18
c1900 n4__i5__bbar vss 159.976e-18
c1901 n16__vdd vss 64.4887e-18
c1902 n14__vdd vss 60.1039e-18
c1903 n4__i3__abar vss 247.657e-18
c1904 n4__i1__net1 vss 79.1509e-18
c1905 n4__i2__net1 vss 62.2602e-18
c1906 n4__i5__abar vss 248.322e-18
c1907 n29__clk4b vss 72.5379e-18
c1908 n3__a0 vss 93.1678e-18
c1909 n16__x0 vss 95.0144e-18
c1910 n13__y0 vss 95.433e-18
c1911 n3__a2 vss 92.5749e-18
c1912 n2__i3__net3 vss 126.859e-18
c1913 n2__i5__net3 vss 139.738e-18
c1914 n6__i3__bbar vss 120.22e-18
c1915 n6__i5__bbar vss 125.506e-18
c1916 n6__i3__abar vss 118.231e-18
c1917 n7__i1__net1 vss 88.6115e-18
c1918 n7__i2__net1 vss 74.0981e-18
c1919 n6__i5__abar vss 112.327e-18
c1920 n131__vdd vss 63.7348e-18
c1921 n36__clk4 vss 32.663e-18
c1922 n12__i0__net4 vss 36.5653e-18
c1923 n6__i0__net3 vss 37.8309e-18
c1924 n7__i0__net6 vss 83.9094e-18
c1925 n33__clk4 vss 50.3984e-18
c1926 n128__vdd vss 55.966e-18
c1927 n14__i0__net4 vss 53.7834e-18
c1928 n130__vdd vss 64.6699e-18
c1929 n7__i0__net3 vss 72.3316e-18
c1930 n133__vdd vss 102.87e-18
c1931 n4__i0__net6 vss 85.4208e-18
c1932 n12__i0__net1 vss 36.5281e-18
c1933 n12__clk2 vss 37.0272e-18
c1934 n8__clkb vss 40.7439e-18
c1935 n7__vdd vss 43.6659e-18
c1936 n7__i0__net2 vss 72.8734e-18
c1937 n14__i0__net1 vss 59.7888e-18
c1938 n136__vdd vss 74.2938e-18
c1939 n11__clk2 vss 47.7007e-18
c1940 n9__clkb vss 87.7939e-18
c1941 n137__vdd vss 158.133e-18
c1942 n5__vdd vss 56.5539e-18
c1943 n4__i0__net2 vss 68.7909e-18
c1944 n4__clk vss 11.8078e-18
c1945 n10__i0__net1 vss 27.8066e-18
c1946 n6__vdd vss 24.6146e-18
c1947 n7__clkb vss 46.7001e-18
c1948 n9__clk2 vss 31.0504e-18
c1949 n10__i0__net4 vss 46.8358e-18
c1950 n5__i0__net3 vss 54.9717e-18
c1951 n13__i0__net4 vss 49.803e-18
c1952 n35__clk4 vss 28.6673e-18
c1953 n5__yin0 vss 50.027e-18
c1954 n10__x2 vss 60.142e-18
c1955 n12__x2 vss 29.1815e-18
c1956 n10__x0 vss 60.4303e-18
c1957 n12__x0 vss 29.4518e-18
c1958 n53__vdd vss 88.2027e-18
c1959 n10__y2 vss 53.3067e-18
c1960 n12__y2 vss 25.4041e-18
c1961 n56__vdd vss 112.723e-18
c1962 n59__vdd vss 107.461e-18
c1963 n2__a2 vss 133.334e-18
c1964 n2__a0 vss 129.862e-18
c1965 n5__yin1 vss 48.9926e-18
c1966 n14__y1 vss 99.5174e-18
c1967 n14__x1 vss 99.2738e-18
c1968 n8__i2__net4 vss 38.2903e-18
c1969 n10__i2__net4 vss 60.5599e-18
c1970 n52__clk4 vss 61.6552e-18
c1971 n53__clk4 vss 47.803e-18
c1972 n55__clk4 vss 62.2326e-18
c1973 n10__i1__rstb vss 70.2948e-18
c1974 n10__x3 vss 58.448e-18
c1975 n5__yin3 vss 41.7365e-18
c1976 n2__c0 vss 53.4825e-18
c1977 n12__y3 vss 24.751e-18
c1978 n21__x1 vss 60.4656e-18
c1979 n75__vdd vss 99.6721e-18
c1980 n47__clk4b vss 227.27e-18
c1981 n48__clk4b vss 262.43e-18
c1982 n51__clk4b vss 264.578e-18
c1983 n52__clk4b vss 215.253e-18
c1984 n62__clk4 vss 115.165e-18
c1985 n63__clk4 vss 166.664e-18
c1986 n65__clk4 vss 139.05e-18
c1987 n67__clk4 vss 115.076e-18
c1988 n2__c1 vss 58.0466e-18
c1989 n37__rst vss 105.428e-18
c1990 n38__rst vss 239.987e-18
c1991 n39__rst vss 149.919e-18
c1992 n40__rst vss 278.479e-18
c1993 n41__rst vss 167.599e-18
c1994 n42__rst vss 112.333e-18
c1995 n2__net12 vss 48.2944e-18
c1996 n97__vdd vss 184.261e-18
c1997 n98__vdd vss 96.8235e-18
c1998 n99__vdd vss 200.988e-18
c1999 n100__vdd vss 172.317e-18
c2000 n101__vdd vss 84.4755e-18
c2001 n102__vdd vss 67.8729e-18
c2002 n112__vdd vss 108.674e-18
c2003 n113__vdd vss 54.2483e-18
c2004 n114__vdd vss 52.4257e-18
c2005 n115__vdd vss 164.841e-18
c2006 n116__vdd vss 148.149e-18
c2007 n117__vdd vss 66.8185e-18
c2008 n118__vdd vss 50.9983e-18
c2009 n126__vdd vss 27.1888e-18
c2010 n127__vdd vss 28.9429e-18
c2011 n129__vdd vss 64.1225e-18
c2012 n132__vdd vss 96.8227e-18
c2013 n134__vdd vss 37.4615e-18
c2014 n135__vdd vss 81.2317e-18
c2015 n22__y1 vss 53.4947e-18
c2016 n24__y1 vss 26.4186e-18
c2017 n6__c0 vss 63.931e-18
c2018 n14__i2__rstb vss 32.958e-18
c2019 n14__i1__rstb vss 32.6872e-18
c2020 n17__i2__rstb vss 445.395e-18
c2021 n17__i1__rstb vss 444.801e-18
c2022 n6__c1 vss 41.8061e-18
c2023 n10__a1 vss 130.794e-18
c2024 n2__i10__net116 vss 58.184e-18
c2025 n10__a3 vss 210.36e-18
c2026 n6__net12 vss 66.2688e-18
c2027 n10__c1 vss 69.03e-18
c2028 n10__c0 vss 45.677e-18
c2029 n10__net12 vss 59.7177e-18
c2030 n14__c1 vss 65.3316e-18
c2031 n14__c0 vss 46.5355e-18
c2032 n7__i8__net51 vss 45.7584e-18
c2033 n7__i7__net51 vss 47.6186e-18
c2034 n11__s1 vss 107.553e-18
c2035 n11__s0 vss 122.556e-18
c2036 n4__i10__net114 vss 17.9199e-18
c2037 n5__i8__carry_bar vss 127.966e-18
c2038 n5__i7__carry_bar vss 131.349e-18
c2039 n153__vdd vss 42.1385e-18
c2040 n154__vdd vss 35.46e-18
c2041 n155__vdd vss 43.8374e-18
c2042 n156__vdd vss 69.5025e-18
c2043 n157__vdd vss 49.3205e-18
c2044 n158__vdd vss 13.2645e-18
c2045 n160__vdd vss 13.5861e-18
c2046 n168__vdd vss 43.2064e-18
c2047 n169__vdd vss 48.5355e-18
c2048 n170__vdd vss 53.6624e-18
c2049 n171__vdd vss 64.5199e-18
c2050 n172__vdd vss 49.9534e-18
c2051 n173__vdd vss 14.8045e-18
c2052 n175__vdd vss 13.6311e-18
c2053 n4__i10__net124 vss 31.413e-18
c2054 n7__i9__net51 vss 47.5052e-18
c2055 n9__i10__net124 vss 26.5903e-18
c2056 n3__r0 vss 89.8411e-18
c2057 n16__i10__net116 vss 10.5758e-18
c2058 n3__i10__net122 vss 26.4697e-18
c2059 n8__i10__net122 vss 26.2387e-18
c2060 n5__i9__carry_bar vss 128.693e-18
c2061 n192__vdd vss 47.7089e-18
c2062 n193__vdd vss 13.25e-18
c2063 n194__vdd vss 52.5591e-18
c2064 n195__vdd vss 104.584e-18
c2065 n196__vdd vss 68.0878e-18
c2066 n197__vdd vss 16.5412e-18
c2067 n199__vdd vss 14.3729e-18
c2068 n2__i14__shift vss 10.4859e-18
c2069 n15__i10__net114 vss 78.041e-18
c2070 n10__i14__shift vss 8.75285e-18
c2071 n208__vdd vss 22.7429e-18
c2072 n209__vdd vss 21.8476e-18
c2073 n210__vdd vss 49.3071e-18
c2074 n211__vdd vss 22.0597e-18
c2075 n212__vdd vss 37.9194e-18
c2076 n213__vdd vss 34.7199e-18
c2077 n214__vdd vss 64.1293e-18
c2078 n215__vdd vss 27.9777e-18
c2079 n2__r2 vss 95.3656e-18
c2080 n18__i14__shift vss 8.64072e-18
c2081 n3__i14__i3__rstb vss 40.5355e-18
c2082 n26__i14__shift vss 49.6484e-18
c2083 n10__i14__i7__net1 vss 47.6235e-18
c2084 n67__rst vss 279.189e-18
c2085 n3__i14__i4__rstb vss 48.1786e-18
c2086 n31__clk vss 658.724e-18
c2087 n32__clk vss 777.139e-18
c2088 n3__i14__i5__rstb vss 48.8901e-18
c2089 n256__vdd vss 99.6887e-18
c2090 n260__vdd vss 65.0341e-18
c2091 n27__clkb vss 226.219e-18
c2092 n28__clkb vss 210.466e-18
c2093 n29__clkb vss 739.799e-18
c2094 n30__clkb vss 771.327e-18
c2095 n39__i14__shift vss 23.3619e-18
c2096 n41__i14__shift vss 24.5177e-18
c2097 n3__vddio vss 29.8754e-18
c2098 n4__i11__net1 vss 33.8667e-18
c2099 n3__net5 vss 76.1143e-18
c2100 n273__vdd vss 11.1583e-18
c2101 n7__r_in vss 56.6782e-18
c2102 n8__r_in vss 137.068e-18
c2103 n8__i12__net1 vss 51.5218e-18
c2104 n11__vddio vss 47.4815e-18
c2105 n12__vddio vss 318.529e-21
c2106 n20__vddio vss 39.2491e-18
c2107 n46__i12__net2 vss 61.5228e-18
c2108 n365__i12__net3 vss 97.1487e-18
c2109 n401__r_out vss 123.697e-18
c2110 n72__rst vss 127.161e-18
c2111 n73__rst vss 71.6815e-18
c2112 n14__serial_out vss 120.873e-18
c2113 n313__vddio vss 107.201e-18
rc1 n314__vddio vddio 425.9e-3
rc3 n165__vss n460__vss 706.6e-3
rc4 n460__vss n461__vss 681.7e-3
rc5 n461__vss n462__vss 527.7e-3
rc7 n129__vss n460__vss 280e-3
rc8 n58__vss n461__vss 280e-3
rc9 n39__vss n462__vss 280e-3
rc11 n465__vss n466__vss 704e-3
rc12 n466__vss n467__vss 683.4e-3
rc13 n467__vss n468__vss 526.8e-3
rc15 n166__vss n465__vss 280e-3
rc16 n127__vss n466__vss 280e-3
rc17 n56__vss n467__vss 280e-3
rc18 n38__vss n468__vss 280e-3
rc19 n457__vss n216__vss 420.3e-3
rc20 n216__vss n168__vss 268.5e-3
rc21 n168__vss n124__vss 234.5e-3
rc22 n124__vss n53__vss 226.6e-3
rc23 n53__vss n36__vss 175.6e-3
rc24 n36__vss n14__vss 231.1e-3
rc25 n457__vss n458__vss 35.08e-3
rc26 n282__vdd n247__vdd 350.6e-3
rc27 n247__vdd n246__vdd 255.5e-3
rc28 n246__vdd n283__vdd 230.5e-3
rc29 n283__vdd n95__vdd 193.7e-3
rc30 n95__vdd n52__vdd 218.4e-3
rc31 n52__vdd n13__vdd 260.3e-3
rc32 n13__vdd vdd 37.95e-3
rc33 n184__vdd n283__vdd 280e-3
rc35 n471__vss n472__vss 705.7e-3
rc36 n472__vss n473__vss 680.9e-3
rc37 n473__vss n474__vss 527.7e-3
rc39 n167__vss n471__vss 280e-3
rc40 n126__vss n472__vss 280e-3
rc41 n55__vss n473__vss 280e-3
rc42 n37__vss n474__vss 280e-3
rd1 n14__vss n13__vss 1.5524
rd2 n13__vdd n12__vdd 545.4e-3
rd3 n36__vss n33__vss 412.3e-3
rd4 n33__vss n37__vss 256.5e-3
rd5 n37__vss n35__vss 137e-3
rd6 n35__vss n38__vss 196e-3
rd7 n38__vss n34__vss 81.32e-3
rd8 n34__vss n39__vss 603.8e-3
rd10 n52__vdd n46__vdd 406.7e-3
rd11 n46__vdd n53__vdd 497.5e-3
rd12 n53__vdd n45__vdd 10.84e-3
rd13 n53__vdd n54__vdd 285.6e-3
rd14 n54__vdd n49__vdd 331.7e-3
rd15 n54__vdd n50__vdd 7.086e-3
rd16 n53__vss n54__vss 393.5e-3
rd17 n54__vss n55__vss 271.9e-3
rd18 n55__vss n56__vss 333.3e-3
rd19 n56__vss n57__vss 505.8e-3
rd20 n57__vss n58__vss 173.7e-3
rd22 n95__vdd n92__vdd 434.6e-3
rd23 n92__vdd n89__vdd 429.8e-3
rd24 n89__vdd n94__vdd 635.7e-3
rd25 n124__vss n125__vss 389.2e-3
rd26 n125__vss n126__vss 277.3e-3
rd27 n126__vss n127__vss 332.7e-3
rd28 n127__vss n128__vss 332.9e-3
rd29 n128__vss n129__vss 349.2e-3
rd31 n140__vdd n183__vdd 1.1522
rd32 n183__vdd n184__vdd 97.09e-3
rd33 n165__vss n163__vss 626.6e-3
rd34 n163__vss n166__vss 328.9e-3
rd35 n166__vss n167__vss 331.8e-3
rd36 n167__vss n164__vss 267.9e-3
rd37 n164__vss n168__vss 390.1e-3
rd38 n243__vdd n246__vdd 429.6e-3
rd39 n243__vdd n244__vdd 855.1e-3
rd40 n215__vss n216__vss 740.5e-3
rd41 n247__vdd n245__vdd 624.1e-3
rd42 n282__vdd n281__vdd 1.5121
rd43 n457__vss n455__vss 591e-3
rd45 n311__vddio n313__vddio 639.6e-3
rd46 n313__vddio n310__vddio 452.1e-3
rd47 n313__vddio n314__vddio 627.8e-3
rd49 n458__vss n456__vss 430.1e-3
re1 n13__vss n12__vss 250e-3
re2 n11__vdd n12__vdd 250e-3
re3 n33__vss n30__vss 250e-3
re4 n34__vss n31__vss 250e-3
re5 n32__vss n35__vss 250e-3
re6 n40__vdd n45__vdd 500e-3
re7 n46__vdd n41__vdd 500e-3
re8 n42__vdd n49__vdd 500e-3
re9 n50__vdd n43__vdd 500e-3
re10 n57__vss n64__vss 500e-3
re11 n65__vss n54__vss 500e-3
re12 n89__vdd n86__vdd 500e-3
re13 n87__vdd n92__vdd 500e-3
re14 n88__vdd n94__vdd 500e-3
re15 n135__vss n128__vss 500e-3
re16 n125__vss n136__vss 500e-3
re18 n143__vdd n183__vdd 250e-3
re19 n161__vss n163__vss 250e-3
re20 n164__vss n162__vss 250e-3
re21 n226__vdd n243__vdd 250e-3
re22 n244__vdd n227__vdd 250e-3
re23 n215__vss n214__vss 250e-3
re24 n242__vdd n245__vdd 250e-3
re25 n310__vddio n308__vddio 250e-3
re26 n281__vdd n280__vdd 250e-3
re27 n453__vss n455__vss 250e-3
re28 n309__vddio n311__vddio 250e-3
re29 n456__vss n454__vss 250e-3
rf1 n12__vss n11__vss 250e-3
rf2 n9__vdd n11__vdd 250e-3
rf3 n30__vss n25__vss 250e-3
rf4 n31__vss n27__vss 250e-3
rf5 n28__vss n32__vss 250e-3
rf17 n140__vdd n141__vdd 500e-3
rf18 n142__vdd n143__vdd 500e-3
rf19 n159__vss n161__vss 250e-3
rf20 n162__vss n160__vss 250e-3
rf21 n224__vdd n226__vdd 250e-3
rf22 n227__vdd n225__vdd 250e-3
rf23 n213__vss n214__vss 250e-3
rf24 n242__vdd n241__vdd 250e-3
rf25 n17__r0 n9__r0 5.6676
rf26 n306__vddio n308__vddio 250e-3
rf27 n279__vdd n280__vdd 250e-3
rf28 n453__vss n451__vss 250e-3
rf29 n309__vddio n307__vddio 250e-3
rf30 n452__vss n454__vss 250e-3
rg1 n3__vss n11__vss 500e-3
rg2 n9__vdd n3__vdd 500e-3
rg3 clk n9__clk 1.8017
rg4 n21__vss n25__vss 500e-3
rg5 n22__vss n27__vss 500e-3
rg6 n28__vss n23__vss 500e-3
rg7 n40__vdd n36__vdd 250e-3
rg8 n37__vdd n41__vdd 250e-3
rg9 n42__vdd n38__vdd 250e-3
rg10 n39__vdd n43__vdd 250e-3
rg11 n62__vss n64__vss 250e-3
rg12 n65__vss n63__vss 250e-3
rg13 n83__vdd n86__vdd 250e-3
rg14 n87__vdd n84__vdd 250e-3
rg15 n88__vdd n85__vdd 250e-3
rg16 n135__vss n133__vss 250e-3
rg17 n134__vss n136__vss 250e-3
rg20 n159__vss n151__vss 250e-3
rg21 n154__vss n160__vss 250e-3
rg22 n224__vdd n205__vdd 250e-3
rg23 n206__vdd n225__vdd 250e-3
rg24 n8__r0 n9__r0 250e-3
rg25 n212__vss n213__vss 250e-3
rg26 n65__rst n67__rst 5.5253
rg27 n67__rst n33__rst 80.29e-3
rg28 n33__rst rst 5.5827
rg29 n67__rst n44__rst 809e-3
rg30 n240__vdd n241__vdd 250e-3
rg31 n17__r0 n16__r0 250e-3
rg32 n304__vddio n306__vddio 250e-3
rg33 n278__vdd n279__vdd 250e-3
rg34 n451__vss n449__vss 250e-3
rg35 n307__vddio n305__vddio 250e-3
rg36 n450__vss n452__vss 250e-3
rh6 n36__vdd n32__vdd 250e-3
rh7 n33__vdd n37__vdd 250e-3
rh8 n38__vdd n34__vdd 250e-3
rh9 n35__vdd n39__vdd 250e-3
rh10 n60__vss n62__vss 250e-3
rh11 n63__vss n61__vss 250e-3
rh12 n80__vdd n83__vdd 250e-3
rh13 n84__vdd n81__vdd 250e-3
rh14 n85__vdd n82__vdd 250e-3
rh15 n32__rst n33__rst 500e-3
rh16 n44__rst n34__rst 500e-3
rh17 n133__vss n131__vss 250e-3
rh18 n132__vss n134__vss 250e-3
rh19 n144__vdd n141__vdd 500e-3
rh20 n142__vdd n147__vdd 500e-3
rh21 n151__vss n152__vss 500e-3
rh22 n153__vss n154__vss 500e-3
rh23 n205__vdd n189__vdd 250e-3
rh24 n190__vdd n206__vdd 250e-3
rh25 n7__r0 n8__r0 500e-3
rh26 n211__vss n212__vss 250e-3
rh27 n65__rst n66__rst 1
rh28 n239__vdd n240__vdd 250e-3
rh30 n31__clk n32__clk 10.9045
rh32 n31__clk n34__clk 2.0672
rh33 n32__clk n9__clk 3.5192
rh35 n12__r1 n7__r1 2.4208
rh36 n15__r0 n16__r0 250e-3
rh37 n304__vddio n302__vddio 250e-3
rh38 n278__vdd n277__vdd 250e-3
rh39 n447__vss n449__vss 250e-3
rh40 n303__vddio n305__vddio 250e-3
rh41 n450__vss n448__vss 250e-3
ri1 n9__clk n10__clk 1
ri2 n2__vss n3__vss 250e-3
ri3 n3__vdd n2__vdd 250e-3
ri4 n11__clkb n10__clkb 2.2977
ri5 n16__vss n21__vss 250e-3
ri6 n18__vss n22__vss 250e-3
ri7 n23__vss n19__vss 250e-3
ri8 n39__clk4b n32__clk4b 1.9793
ri9 n23__vdd n32__vdd 250e-3
ri10 n33__vdd n24__vdd 250e-3
ri11 n27__vdd n34__vdd 250e-3
ri12 n35__vdd n28__vdd 250e-3
ri13 n14__y0 n15__y0 2.0362
ri14 n18__x0 n19__x0 2.3158
ri15 n17__x0 n19__x0 500e-3
ri16 n60__vss n49__vss 250e-3
ri17 n52__vss n61__vss 250e-3
ri18 n18__y1 n6__y1 737.1e-3
ri19 n18__x1 n10__x1 737.1e-3
ri20 n18__x2 n14__x2 2.8531
ri21 n18__y2 n14__y2 3.7804
ri22 n24__x1 n12__x1 3.0228
ri23 n80__vdd n67__vdd 250e-3
ri24 n69__vdd n81__vdd 250e-3
ri25 n77__vdd n82__vdd 250e-3
ri26 n21__y1 n12__y1 2.4681
ri27 n15__y3 n13__y3 3.0639
ri28 n14__x3 n13__x3 2.5166
ri29 n31__rst n32__rst 1
ri30 n34__rst n35__rst 1
ri31 n131__vss n120__vss 250e-3
ri32 n123__vss n132__vss 250e-3
ri35 n15__s1 n14__s1 4.1101
ri36 n152__vss n155__vss 250e-3
ri37 n156__vss n153__vss 250e-3
ri38 n189__vdd n185__vdd 250e-3
ri39 n188__vdd n190__vdd 250e-3
ri40 n7__r0 n6__r0 1.4621
ri41 n7__r1 n4__r1 1
ri42 n210__vss n211__vss 250e-3
ri43 n74__clk4 n66__clk4 9.4305
ri44 n22__clk2 n13__clk2 11.7382
ri45 n235__vdd n239__vdd 250e-3
ri46 n237__vdd n238__vdd 618.5e-3
ri47 n220__vss n222__vss 464.4e-3
ri48 n4__i14__net2 n5__i14__net2 1.4421
ri49 n9__r2 n5__r2 2.3357
ri50 n10__i14__net9 n6__i14__net9 1.2289
ri51 n8__i14__net8 n9__i14__net8 480.8e-3
ri52 n71__rst n72__rst 888.1e-3
ri53 n72__rst n73__rst 828.4e-3
ri54 n73__rst n66__rst 419e-3
ri55 n72__rst n69__rst 30.6e-3
ri56 n73__rst n64__rst 51.3e-3
ri57 n11__r1 n12__r1 500e-3
ri58 n10__i14__net15 n6__i14__net15 1.3659
ri59 n7__i14__net14 n9__i14__net14 434.9e-3
ri60 n14__r0 n15__r0 250e-3
ri61 n39__clk n41__clk 1.3499
ri62 n41__clk n34__clk 618.8e-3
ri63 n34__clk n28__clk 720.1e-3
ri64 n36__clk n41__clk 500e-3
ri65 n13__serial_out n14__serial_out 1.0961
ri67 n14__serial_out n11__serial_out 273.6e-3
ri68 n7__vddio n302__vddio 250e-3
ri69 n277__vdd n269__vdd 250e-3
ri70 n251__vss n447__vss 250e-3
ri71 n9__vddio n303__vddio 250e-3
ri72 n448__vss n255__vss 250e-3
rj1 n1__vss n2__vss 500e-3
rj2 n1__vdd n2__vdd 500e-3
rj3 n9__i0__net2 n6__i0__net2 824.8e-3
rj4 n13__clk n11__clk 810.9e-3
rj5 n11__clk n12__clk 1.3804
rj6 n12__clk n10__clk 208.3e-3
rj7 n6__clkb n10__clkb 250e-3
rj8 n11__i0__net1 n9__i0__net1 1.5922
rj9 n16__i0__net1 n13__i0__net1 1.3296
rj10 n9__i0__net6 n6__i0__net6 825.1e-3
rj11 n15__clk2 n14__clk2 806.8e-3
rj12 n14__clk2 n13__clk2 213.1e-3
rj14 n13__clk2 n10__clk2 830.2e-3
rj15 n11__i0__net4 n9__i0__net4 1.5949
rj16 n15__vss n16__vss 500e-3
rj17 n17__vss n18__vss 500e-3
rj18 n19__vss n20__vss 500e-3
rj19 n22__vdd n23__vdd 500e-3
rj20 n24__vdd n25__vdd 500e-3
rj21 n26__vdd n27__vdd 500e-3
rj22 n28__vdd n29__vdd 500e-3
rj23 n30__vdd n19__vdd 710.4e-3
rj24 n19__vdd n15__vdd 213.5e-3
rj25 n11__x2 n13__x2 797.2e-3
rj26 n13__x2 n14__x2 501.9e-3
rj27 n8__x2 n13__x2 500e-3
rj28 n31__vdd n21__vdd 710.4e-3
rj29 n21__vdd n17__vdd 213.5e-3
rj30 n11__x0 n17__x0 794.8e-3
rj31 n17__x0 n8__x0 501.9e-3
rj32 n10__y0 n14__y0 1
rj33 n18__x0 n13__x0 1
rj34 n5__y1 n6__y1 500e-3
rj35 n10__x1 n9__x1 500e-3
rj36 n45__vss n48__vss 1.0132
rj37 n11__y2 n13__y2 973.9e-3
rj38 n13__y2 n14__y2 501.9e-3
rj39 n9__y2 n13__y2 500e-3
rj40 n47__vss n42__vss 1.0132
rj41 n10__i2__net1 n11__i2__net1 345.5e-3
rj42 n11__i2__net1 n6__i2__net1 299.6e-3
rj43 n8__i2__net1 n11__i2__net1 500e-3
rj44 n10__i1__net1 n11__i1__net1 345.5e-3
rj45 n11__i1__net1 n6__i1__net1 299.6e-3
rj46 n8__i1__net1 n11__i1__net1 500e-3
rj47 n17__y0 n19__y0 969e-3
rj48 n19__y0 n15__y0 1.802e-3
rj49 n9__y0 n19__y0 500e-3
rj50 n49__vss n50__vss 500e-3
rj51 n51__vss n52__vss 500e-3
rj52 n6__i2__net3 n8__i2__net3 802.2e-3
rj53 n6__i1__net3 n8__i1__net3 802.2e-3
rj54 n11__y1 n12__y1 1.0634
rj55 n11__x1 n12__x1 1.0634
rj56 n13__y1 n18__y1 503.6e-3
rj57 n13__x1 n18__x1 503.6e-3
rj58 n16__y2 n18__y2 1
rj59 n18__x2 n16__x2 1
rj60 n65__vdd n64__vdd 710.4e-3
rj61 n64__vdd n62__vdd 213.5e-3
rj62 n11__x3 n13__x3 795.5e-3
rj63 n13__x3 n8__x3 500e-3
rj64 n66__vdd n67__vdd 500e-3
rj65 n68__vdd n69__vdd 500e-3
rj66 n77__vdd n78__vdd 500e-3
rj67 n45__clk4b n47__clk4b 1.2275
rj68 n47__clk4b n48__clk4b 561.6e-3
rj69 n48__clk4b n39__clk4b 950.9e-3
rj71 n47__clk4b n43__clk4b 555.2e-3
rj72 n48__clk4b n41__clk4b 555.2e-3
rj73 n37__clk4b n39__clk4b 500e-3
rj75 n32__clk4b n50__clk4b 394.4e-3
rj76 n50__clk4b n51__clk4b 948.4e-3
rj77 n51__clk4b n42__clk4b 555.2e-3
rj78 n51__clk4b n52__clk4b 561.6e-3
rj79 n52__clk4b n44__clk4b 555.2e-3
rj80 n52__clk4b n46__clk4b 1.2272
rj81 n38__clk4b n50__clk4b 500e-3
rj82 n78__vss n71__vss 1.0132
rj83 n11__y3 n13__y3 958e-3
rj84 n13__y3 n9__y3 512.1e-3
rj85 n6__i2__net2 n8__i2__net2 832.7e-3
rj86 n6__i1__net2 n8__i1__net2 832.7e-3
rj87 n79__vdd n73__vdd 710.4e-3
rj88 n73__vdd n71__vdd 213.5e-3
rj89 n60__clk4 n58__clk4 843.7e-3
rj90 n58__clk4 n61__clk4 511.4e-3
rj91 n61__clk4 n50__clk4 348.5e-3
rj92 n50__clk4 n62__clk4 329.6e-3
rj93 n62__clk4 n48__clk4 569.7e-3
rj94 n62__clk4 n46__clk4 270.2e-3
rj95 n46__clk4 n63__clk4 784.1e-3
rj96 n63__clk4 n44__clk4 569.7e-3
rj97 n63__clk4 n42__clk4 247.6e-3
rj98 n42__clk4 n64__clk4 440.6e-3
rj99 n64__clk4 n41__clk4 1.1678
rj100 n41__clk4 n65__clk4 244e-3
rj101 n65__clk4 n43__clk4 569.7e-3
rj102 n64__clk4 n66__clk4 990.7e-3
rj103 n65__clk4 n45__clk4 783.9e-3
rj104 n45__clk4 n67__clk4 270.2e-3
rj105 n67__clk4 n47__clk4 569.7e-3
rj106 n67__clk4 n49__clk4 329.6e-3
rj107 n49__clk4 n68__clk4 348.4e-3
rj108 n68__clk4 n57__clk4 511e-3
rj109 n57__clk4 n59__clk4 843.3e-3
rj110 n54__clk4 n61__clk4 500e-3
rj111 n34__clk4 n64__clk4 500e-3
rj112 n51__clk4 n68__clk4 500e-3
rj113 n22__x1 n24__x1 793.5e-3
rj114 n24__x1 n19__x1 500e-3
rj115 n14__y3 n15__y3 1
rj116 n14__x3 n15__x3 1
rj117 n11__i2__net4 n12__i2__net4 1.5661
rj118 n12__i2__net4 n6__i2__net4 302e-3
rj119 n9__i2__net4 n12__i2__net4 500e-3
rj120 n11__i1__net4 n12__i1__net4 1.5661
rj121 n12__i1__net4 n6__i1__net4 302e-3
rj122 n9__i1__net4 n12__i1__net4 500e-3
rj123 n36__rst n37__rst 825.7e-3
rj124 n37__rst n38__rst 630.6e-3
rj125 n38__rst n39__rst 1.2252
rj126 n39__rst n17__rst 679.8e-3
rj127 n37__rst n31__rst 125.3e-3
rj128 n38__rst n29__rst 515.2e-3
rj129 n39__rst n19__rst 515.2e-3
rj130 n30__rst n40__rst 515.2e-3
rj131 n40__rst n41__rst 1.2252
rj132 n41__rst n18__rst 679.8e-3
rj133 n40__rst n42__rst 695.1e-3
rj134 n42__rst n35__rst 90.16e-3
rj135 n41__rst n20__rst 515.2e-3
rj136 n42__rst n43__rst 727.1e-3
rj137 n15__i2__rstb n17__i2__rstb 840e-3
rj138 n17__i2__rstb n9__i2__rstb 1.7949
rj139 n17__i2__rstb n11__i2__rstb 550.4e-3
rj140 n15__i1__rstb n17__i1__rstb 840e-3
rj141 n17__i1__rstb n9__i1__rstb 1.7949
rj142 n17__i1__rstb n11__i1__rstb 550.4e-3
rj143 n119__vss n75__vss 1.0132
rj144 n23__y1 n21__y1 973.6e-3
rj145 n21__y1 n20__y1 500e-3
rj146 n120__vss n121__vss 500e-3
rj147 n122__vss n123__vss 500e-3
rj148 n148__vdd n144__vdd 500e-3
rj149 n147__vdd n151__vdd 500e-3
rj150 n4__i8__net51 n9__i8__net51 1.3312
rj151 n4__i7__net51 n9__i7__net51 1.3285
rj152 n10__s1 n14__s1 1
rj153 n17__a2 n18__a2 904.4e-3
rj154 n18__a2 n4__a2 3.7738
rj155 n16__a2 n17__a2 500e-3
rj156 n13__a2 n18__a2 500e-3
rj157 n17__a0 n18__a0 853e-3
rj158 n18__a0 n4__a0 3.1864
rj159 n16__a0 n17__a0 500e-3
rj160 n13__a0 n18__a0 500e-3
rj161 n9__a3 n13__a3 653.3e-3
rj162 n13__a3 n14__a3 800.4e-3
rj163 n15__a1 n13__a1 1.3925
rj164 n13__a1 n12__a1 1.3377
rj165 n19__c0 n21__c0 1.4267
rj166 n18__c1 n20__c1 1.5961
rj167 n9__i10__net116 n10__i10__net116 1.3624
rj168 n155__vss n157__vss 250e-3
rj169 n158__vss n156__vss 250e-3
rj170 n4__i9__net51 n9__i9__net51 1.3419
rj171 i10__net115 n2__i10__net115 1.1542
rj172 i10__net124 n2__i10__net124 1.1581
rj173 n2__r0 n6__r0 1
rj174 n17__net12 n15__net12 3.3403
rj175 n18__s0 n19__s0 890.2e-3
rj176 n19__s0 n10__s0 1.6239
rj177 n17__s0 n18__s0 500e-3
rj178 n14__s0 n19__s0 500e-3
rj179 n4__i10__net125 i10__net125 1.1581
rj180 i10__net122 n4__i10__net122 1.1619
rj181 n185__vdd n186__vdd 500e-3
rj182 n187__vdd n188__vdd 500e-3
rj183 n18__s1 n16__s1 1.3459
rj184 n16__s1 n15__s1 19.82e-3
rj185 n12__i10__net114 n15__i10__net114 85.23e-3
rj186 n15__i10__net114 n8__i10__net114 416.2e-3
rj187 n15__i10__net114 n16__i10__net114 900.7e-3
rj188 n17__i10__net114 n14__i10__net114 927e-3
rj189 n14__i10__net114 n9__i10__net114 443.7e-3
rj190 n18__i10__net116 n19__i10__net116 2.1819
rj192 n4__r1 n5__r1 75.17e-3
rj193 n5__r1 n2__r1 763.1e-3
rj194 n5__r2 r2 250e-3
rj195 n209__vss n210__vss 500e-3
rj196 n72__clk4 n74__clk4 3.3509
rj197 n20__clk2 n22__clk2 3.64
rj198 n63__rst n64__rst 1.2271
rj199 n9__i14__i7__net1 n10__i14__i7__net1 122.4e-3
rj200 n10__i14__i7__net1 n6__i14__i7__net1 222.6e-3
rj201 n10__i14__i7__net1 n8__i14__i7__net1 167.3e-3
rj202 n234__vdd n235__vdd 500e-3
rj203 n236__vdd n237__vdd 1.3044
rj204 n238__vdd n231__vdd 1.1406
rj205 n28__clk n29__clk 2.416e-3
rj206 n29__clk n27__clk 815.3e-3
rj207 n9__i14__i3__net5 n5__i14__i3__net5 825.9e-3
rj208 n6__i14__net9 n2__i14__net9 2.072
rj209 n248__vdd n232__vdd 1.3839
rj210 n51__rst n69__rst 1.2295
rj211 n220__vss n218__vss 1
rj212 n221__vss n222__vss 1
rj213 n6__i14__i0__net1 n5__i14__i0__net1 886.2e-3
rj214 n4__i14__net2 n6__i14__net2 500e-3
rj215 n5__i14__net2 n7__i14__net2 710.7e-3
rj216 n7__r2 n9__r2 1
rj217 n6__i14__net15 n2__i14__net15 1.6392
rj218 n10__i14__net9 n8__i14__net9 1
rj220 n36__clk n35__clk 815.3e-3
rj221 n8__i14__i1__net1 n5__i14__i1__net1 887e-3
rj222 n9__i14__i4__net5 n5__i14__i4__net5 825.9e-3
rj223 n8__i14__net8 n6__i14__net8 1
rj224 n9__i14__net8 n4__i14__net8 802.9e-3
rj225 n265__vdd n251__vdd 1.3954
rj226 n70__rst n71__rst 1.2295
rj227 n9__r1 n11__r1 1.6721
rj228 n7__serial_out n11__serial_out 1
rj229 n10__i14__net15 n8__i14__net15 1
rj230 n6__i14__i2__net1 n5__i14__i2__net1 887e-3
rj231 n7__i14__net14 n5__i14__net14 1
rj232 n8__i14__net14 n9__i14__net14 1.2614
rj233 n26__clkb n27__clkb 1.6654
rj234 n27__clkb n28__clkb 866e-3
rj235 n28__clkb n29__clkb 1.134
rj236 n29__clkb n30__clkb 12.6653
rj237 n30__clkb n11__clkb 196.8e-3
rj238 n27__clkb n25__clkb 806e-3
rj239 n28__clkb n24__clkb 864.4e-3
rj241 n30__clkb clkb 788.1e-3
rj242 n37__i14__shift n38__i14__shift 693.2e-3
rj243 n38__i14__shift n35__i14__shift 245.4e-3
rj244 n35__i14__shift n39__i14__shift 155.2e-3
rj245 n39__i14__shift n40__i14__shift 149.4e-3
rj246 n40__i14__shift n32__i14__shift 245.4e-3
rj247 n32__i14__shift n41__i14__shift 158.3e-3
rj248 n41__i14__shift n42__i14__shift 149.4e-3
rj249 n42__i14__shift n29__i14__shift 249.2e-3
rj250 n29__i14__shift n25__i14__shift 509.2e-3
rj251 n39__i14__shift n34__i14__shift 540.3e-3
rj252 n41__i14__shift n31__i14__shift 540.3e-3
rj253 n36__i14__shift n38__i14__shift 500e-3
rj254 n33__i14__shift n40__i14__shift 500e-3
rj255 n30__i14__shift n42__i14__shift 500e-3
rj256 n13__r0 n14__r0 250e-3
rj258 n39__clk n38__clk 815.4e-3
rj259 n9__i14__i5__net5 n5__i14__i5__net5 797.2e-3
rj260 n13__serial_out n12__serial_out 1
rj261 n6__vddio n7__vddio 250e-3
rj262 n7__i11__net1 n5__i11__net1 732.2e-3
rj263 n269__vdd n270__vdd 500e-3
rj264 n250__vss n251__vss 500e-3
rj265 n8__vddio n9__vddio 500e-3
rj266 n255__vss n256__vss 500e-3
rj267 n41__i12__net2 n34__i12__net2 1.3247
rj268 n42__i12__net2 n37__i12__net2 1.2616
rj269 n45__vddio n46__vddio 824.7e-3
rj270 n46__vddio n47__vddio 332e-3
rj271 n47__vddio n48__vddio 329.6e-3
rj272 n48__vddio n49__vddio 327.1e-3
rj273 n49__vddio n19__vddio 829.6e-3
rj274 n41__vddio n46__vddio 500e-3
rj275 n37__vddio n47__vddio 500e-3
rj276 n33__vddio n48__vddio 500e-3
rj277 n29__vddio n49__vddio 500e-3
rj278 n290__vss n291__vss 824.7e-3
rj279 n291__vss n292__vss 332e-3
rj280 n292__vss n293__vss 329.6e-3
rj281 n293__vss n294__vss 327.1e-3
rj282 n294__vss n260__vss 829.6e-3
rj283 n286__vss n291__vss 500e-3
rj284 n282__vss n292__vss 500e-3
rj285 n278__vss n293__vss 500e-3
rj286 n274__vss n294__vss 500e-3
rj287 n90__i12__net3 n91__i12__net3 824.7e-3
rj288 n91__i12__net3 n92__i12__net3 334.2e-3
rj289 n92__i12__net3 n93__i12__net3 331.8e-3
rj290 n93__i12__net3 n94__i12__net3 329.3e-3
rj291 n94__i12__net3 n14__i12__net3 831.8e-3
rj292 n78__i12__net3 n91__i12__net3 500e-3
rj293 n62__i12__net3 n92__i12__net3 500e-3
rj294 n46__i12__net3 n93__i12__net3 500e-3
rj295 n30__i12__net3 n94__i12__net3 500e-3
rj296 n95__i12__net3 n96__i12__net3 826.9e-3
rj297 n96__i12__net3 n97__i12__net3 334.2e-3
rj298 n97__i12__net3 n98__i12__net3 331.8e-3
rj299 n98__i12__net3 n99__i12__net3 329.3e-3
rj300 n99__i12__net3 n17__i12__net3 831.8e-3
rj301 n81__i12__net3 n96__i12__net3 500e-3
rj302 n65__i12__net3 n97__i12__net3 500e-3
rj303 n49__i12__net3 n98__i12__net3 500e-3
rj304 n33__i12__net3 n99__i12__net3 500e-3
rj305 n407__r_out n410__r_out 827.1e-3
rj306 n410__r_out n411__r_out 327.1e-3
rj307 n411__r_out n412__r_out 334.4e-3
rj308 n412__r_out n413__r_out 327.1e-3
rj309 n413__r_out n414__r_out 327.1e-3
rj310 n414__r_out n415__r_out 334.4e-3
rj311 n415__r_out n416__r_out 327.1e-3
rj312 n416__r_out n417__r_out 327.1e-3
rj313 n417__r_out n418__r_out 334.4e-3
rj314 n418__r_out n419__r_out 327.1e-3
rj315 n419__r_out n420__r_out 327.1e-3
rj316 n420__r_out n421__r_out 327.1e-3
rj317 n421__r_out n422__r_out 327.1e-3
rj318 n422__r_out n423__r_out 327.1e-3
rj319 n423__r_out n424__r_out 334.4e-3
rj320 n424__r_out n425__r_out 327.1e-3
rj321 n425__r_out n426__r_out 327.1e-3
rj322 n426__r_out n427__r_out 334.4e-3
rj323 n427__r_out n428__r_out 327.1e-3
rj324 n428__r_out n429__r_out 327.1e-3
rj325 n429__r_out n430__r_out 334.4e-3
rj326 n430__r_out n431__r_out 327.1e-3
rj327 n431__r_out n432__r_out 327.1e-3
rj328 n432__r_out n433__r_out 341.6e-3
rj329 n433__r_out n434__r_out 327.1e-3
rj330 n434__r_out n435__r_out 334.4e-3
rj331 n435__r_out n436__r_out 327.1e-3
rj332 n436__r_out n437__r_out 322.3e-3
rj333 n437__r_out n438__r_out 339.2e-3
rj334 n438__r_out n439__r_out 327.1e-3
rj335 n439__r_out n440__r_out 327.1e-3
rj336 n440__r_out n441__r_out 334.4e-3
rj337 n441__r_out n442__r_out 327.1e-3
rj338 n442__r_out n443__r_out 327.1e-3
rj339 n443__r_out n444__r_out 327.1e-3
rj340 n444__r_out n445__r_out 327.1e-3
rj341 n445__r_out n446__r_out 327.1e-3
rj342 n446__r_out n447__r_out 334.4e-3
rj343 n447__r_out n448__r_out 327.1e-3
rj344 n448__r_out n449__r_out 327.1e-3
rj345 n449__r_out n450__r_out 339.2e-3
rj346 n450__r_out n451__r_out 327.1e-3
rj347 n451__r_out n452__r_out 327.1e-3
rj348 n452__r_out n453__r_out 334.4e-3
rj349 n453__r_out n454__r_out 327.1e-3
rj350 n454__r_out n455__r_out 327.1e-3
rj351 n455__r_out n456__r_out 332e-3
rj352 n456__r_out n457__r_out 334.4e-3
rj353 n457__r_out n458__r_out 327.1e-3
rj354 n458__r_out n4__r_out 827.1e-3
rj355 n396__r_out n410__r_out 500e-3
rj356 n388__r_out n411__r_out 500e-3
rj357 n380__r_out n412__r_out 500e-3
rj358 n372__r_out n413__r_out 500e-3
rj359 n364__r_out n414__r_out 500e-3
rj360 n356__r_out n415__r_out 500e-3
rj361 n348__r_out n416__r_out 500e-3
rj362 n340__r_out n417__r_out 500e-3
rj363 n332__r_out n418__r_out 500e-3
rj364 n324__r_out n419__r_out 500e-3
rj365 n316__r_out n420__r_out 500e-3
rj366 n308__r_out n421__r_out 500e-3
rj367 n300__r_out n422__r_out 500e-3
rj368 n292__r_out n423__r_out 500e-3
rj369 n284__r_out n424__r_out 500e-3
rj370 n276__r_out n425__r_out 500e-3
rj371 n268__r_out n426__r_out 500e-3
rj372 n260__r_out n427__r_out 500e-3
rj373 n252__r_out n428__r_out 500e-3
rj374 n244__r_out n429__r_out 500e-3
rj375 n236__r_out n430__r_out 500e-3
rj376 n228__r_out n431__r_out 500e-3
rj377 n220__r_out n432__r_out 500e-3
rj378 n212__r_out n433__r_out 500e-3
rj379 n204__r_out n434__r_out 500e-3
rj380 n196__r_out n435__r_out 500e-3
rj381 n188__r_out n436__r_out 500e-3
rj382 n184__r_out n437__r_out 500e-3
rj383 n172__r_out n438__r_out 500e-3
rj384 n164__r_out n439__r_out 500e-3
rj385 n156__r_out n440__r_out 500e-3
rj386 n148__r_out n441__r_out 500e-3
rj387 n140__r_out n442__r_out 500e-3
rj388 n132__r_out n443__r_out 500e-3
rj389 n124__r_out n444__r_out 500e-3
rj390 n116__r_out n445__r_out 500e-3
rj391 n108__r_out n446__r_out 500e-3
rj392 n100__r_out n447__r_out 500e-3
rj393 n92__r_out n448__r_out 500e-3
rj394 n84__r_out n449__r_out 500e-3
rj395 n76__r_out n450__r_out 500e-3
rj396 n68__r_out n451__r_out 500e-3
rj397 n60__r_out n452__r_out 500e-3
rj398 n52__r_out n453__r_out 500e-3
rj399 n44__r_out n454__r_out 500e-3
rj400 n36__r_out n455__r_out 500e-3
rj401 n28__r_out n456__r_out 500e-3
rj402 n20__r_out n457__r_out 500e-3
rj403 n12__r_out n458__r_out 500e-3
rj404 n402__r_out n459__r_out 827.1e-3
rj405 n459__r_out n460__r_out 327.1e-3
rj406 n460__r_out n461__r_out 334.4e-3
rj407 n461__r_out n462__r_out 327.1e-3
rj408 n462__r_out n463__r_out 327.1e-3
rj409 n463__r_out n464__r_out 334.4e-3
rj410 n464__r_out n465__r_out 327.1e-3
rj411 n465__r_out n466__r_out 327.1e-3
rj412 n466__r_out n467__r_out 334.4e-3
rj413 n467__r_out n468__r_out 327.1e-3
rj414 n468__r_out n469__r_out 327.1e-3
rj415 n469__r_out n470__r_out 327.1e-3
rj416 n470__r_out n471__r_out 327.1e-3
rj417 n471__r_out n472__r_out 327.1e-3
rj418 n472__r_out n473__r_out 334.4e-3
rj419 n473__r_out n474__r_out 327.1e-3
rj420 n474__r_out n475__r_out 327.1e-3
rj421 n475__r_out n476__r_out 334.4e-3
rj422 n476__r_out n477__r_out 327.1e-3
rj423 n477__r_out n478__r_out 327.1e-3
rj424 n478__r_out n479__r_out 334.4e-3
rj425 n479__r_out n480__r_out 327.1e-3
rj426 n480__r_out n481__r_out 327.1e-3
rj427 n481__r_out n482__r_out 341.6e-3
rj428 n482__r_out n483__r_out 327.1e-3
rj429 n483__r_out n484__r_out 334.4e-3
rj430 n484__r_out n485__r_out 327.1e-3
rj431 n485__r_out n486__r_out 327.1e-3
rj432 n486__r_out n487__r_out 334.4e-3
rj433 n487__r_out n488__r_out 327.1e-3
rj434 n488__r_out n489__r_out 327.1e-3
rj435 n489__r_out n490__r_out 334.4e-3
rj436 n490__r_out n491__r_out 327.1e-3
rj437 n491__r_out n492__r_out 327.1e-3
rj438 n492__r_out n493__r_out 327.1e-3
rj439 n493__r_out n494__r_out 327.1e-3
rj440 n494__r_out n495__r_out 327.1e-3
rj441 n495__r_out n496__r_out 334.4e-3
rj442 n496__r_out n497__r_out 327.1e-3
rj443 n497__r_out n498__r_out 327.1e-3
rj444 n498__r_out n499__r_out 339.2e-3
rj445 n499__r_out n500__r_out 327.1e-3
rj446 n500__r_out n501__r_out 327.1e-3
rj447 n501__r_out n502__r_out 334.4e-3
rj448 n502__r_out n503__r_out 327.1e-3
rj449 n503__r_out n504__r_out 327.1e-3
rj450 n504__r_out n505__r_out 332e-3
rj451 n505__r_out n506__r_out 334.4e-3
rj452 n506__r_out n507__r_out 327.1e-3
rj453 n507__r_out n6__r_out 827.1e-3
rj454 n398__r_out n459__r_out 500e-3
rj455 n390__r_out n460__r_out 500e-3
rj456 n382__r_out n461__r_out 500e-3
rj457 n374__r_out n462__r_out 500e-3
rj458 n366__r_out n463__r_out 500e-3
rj459 n358__r_out n464__r_out 500e-3
rj460 n350__r_out n465__r_out 500e-3
rj461 n342__r_out n466__r_out 500e-3
rj462 n334__r_out n467__r_out 500e-3
rj463 n326__r_out n468__r_out 500e-3
rj464 n318__r_out n469__r_out 500e-3
rj465 n310__r_out n470__r_out 500e-3
rj466 n302__r_out n471__r_out 500e-3
rj467 n294__r_out n472__r_out 500e-3
rj468 n286__r_out n473__r_out 500e-3
rj469 n278__r_out n474__r_out 500e-3
rj470 n270__r_out n475__r_out 500e-3
rj471 n262__r_out n476__r_out 500e-3
rj472 n254__r_out n477__r_out 500e-3
rj473 n246__r_out n478__r_out 500e-3
rj474 n238__r_out n479__r_out 500e-3
rj475 n230__r_out n480__r_out 500e-3
rj476 n222__r_out n481__r_out 500e-3
rj477 n214__r_out n482__r_out 500e-3
rj478 n206__r_out n483__r_out 500e-3
rj479 n198__r_out n484__r_out 500e-3
rj480 n190__r_out n485__r_out 500e-3
rj481 n178__r_out n486__r_out 500e-3
rj482 n174__r_out n487__r_out 500e-3
rj483 n166__r_out n488__r_out 500e-3
rj484 n158__r_out n489__r_out 500e-3
rj485 n150__r_out n490__r_out 500e-3
rj486 n142__r_out n491__r_out 500e-3
rj487 n134__r_out n492__r_out 500e-3
rj488 n126__r_out n493__r_out 500e-3
rj489 n118__r_out n494__r_out 500e-3
rj490 n110__r_out n495__r_out 500e-3
rj491 n102__r_out n496__r_out 500e-3
rj492 n94__r_out n497__r_out 500e-3
rj493 n86__r_out n498__r_out 500e-3
rj494 n78__r_out n499__r_out 500e-3
rj495 n70__r_out n500__r_out 500e-3
rj496 n62__r_out n501__r_out 500e-3
rj497 n54__r_out n502__r_out 500e-3
rj498 n46__r_out n503__r_out 500e-3
rj499 n38__r_out n504__r_out 500e-3
rj500 n30__r_out n505__r_out 500e-3
rj501 n22__r_out n506__r_out 500e-3
rj502 n14__r_out n507__r_out 500e-3
rj503 n251__vddio n252__vddio 399.6e-3
rj504 n252__vddio n253__vddio 327.1e-3
rj505 n253__vddio n254__vddio 334.4e-3
rj506 n254__vddio n255__vddio 327.1e-3
rj507 n255__vddio n256__vddio 327.1e-3
rj508 n256__vddio n257__vddio 334.4e-3
rj509 n257__vddio n258__vddio 327.1e-3
rj510 n258__vddio n259__vddio 327.1e-3
rj511 n259__vddio n260__vddio 334.4e-3
rj512 n260__vddio n261__vddio 327.1e-3
rj513 n261__vddio n262__vddio 327.1e-3
rj514 n262__vddio n263__vddio 327.1e-3
rj515 n263__vddio n264__vddio 327.1e-3
rj516 n264__vddio n265__vddio 327.1e-3
rj517 n265__vddio n266__vddio 334.4e-3
rj518 n266__vddio n267__vddio 327.1e-3
rj519 n267__vddio n268__vddio 327.1e-3
rj520 n268__vddio n269__vddio 334.4e-3
rj521 n269__vddio n270__vddio 327.1e-3
rj522 n270__vddio n271__vddio 327.1e-3
rj523 n271__vddio n272__vddio 334.4e-3
rj524 n272__vddio n273__vddio 327.1e-3
rj525 n273__vddio n274__vddio 327.1e-3
rj526 n274__vddio n275__vddio 341.6e-3
rj527 n275__vddio n276__vddio 327.1e-3
rj528 n276__vddio n277__vddio 334.4e-3
rj529 n277__vddio n278__vddio 327.1e-3
rj530 n278__vddio n279__vddio 327.1e-3
rj531 n279__vddio n280__vddio 334.4e-3
rj532 n280__vddio n281__vddio 327.1e-3
rj533 n281__vddio n282__vddio 327.1e-3
rj534 n282__vddio n283__vddio 334.4e-3
rj535 n283__vddio n284__vddio 327.1e-3
rj536 n284__vddio n285__vddio 327.1e-3
rj537 n285__vddio n286__vddio 327.1e-3
rj538 n286__vddio n287__vddio 327.1e-3
rj539 n287__vddio n288__vddio 327.1e-3
rj540 n288__vddio n289__vddio 334.4e-3
rj541 n289__vddio n290__vddio 327.1e-3
rj542 n290__vddio n291__vddio 327.1e-3
rj543 n291__vddio n292__vddio 339.2e-3
rj544 n292__vddio n293__vddio 327.1e-3
rj545 n293__vddio n294__vddio 327.1e-3
rj546 n294__vddio n295__vddio 334.4e-3
rj547 n295__vddio n296__vddio 327.1e-3
rj548 n296__vddio n297__vddio 327.1e-3
rj549 n297__vddio n298__vddio 332e-3
rj550 n298__vddio n299__vddio 334.4e-3
rj551 n299__vddio n300__vddio 327.1e-3
rj552 n300__vddio n301__vddio 331.3e-3
rj553 n301__vddio n24__vddio 4.9414
rj554 n249__vddio n252__vddio 500e-3
rj555 n245__vddio n253__vddio 500e-3
rj556 n241__vddio n254__vddio 500e-3
rj557 n237__vddio n255__vddio 500e-3
rj558 n233__vddio n256__vddio 500e-3
rj559 n229__vddio n257__vddio 500e-3
rj560 n225__vddio n258__vddio 500e-3
rj561 n221__vddio n259__vddio 500e-3
rj562 n217__vddio n260__vddio 500e-3
rj563 n213__vddio n261__vddio 500e-3
rj564 n209__vddio n262__vddio 500e-3
rj565 n205__vddio n263__vddio 500e-3
rj566 n201__vddio n264__vddio 500e-3
rj567 n197__vddio n265__vddio 500e-3
rj568 n193__vddio n266__vddio 500e-3
rj569 n189__vddio n267__vddio 500e-3
rj570 n185__vddio n268__vddio 500e-3
rj571 n181__vddio n269__vddio 500e-3
rj572 n177__vddio n270__vddio 500e-3
rj573 n173__vddio n271__vddio 500e-3
rj574 n169__vddio n272__vddio 500e-3
rj575 n165__vddio n273__vddio 500e-3
rj576 n161__vddio n274__vddio 500e-3
rj577 n157__vddio n275__vddio 500e-3
rj578 n153__vddio n276__vddio 500e-3
rj579 n149__vddio n277__vddio 500e-3
rj580 n145__vddio n278__vddio 500e-3
rj581 n141__vddio n279__vddio 500e-3
rj582 n136__vddio n280__vddio 500e-3
rj583 n132__vddio n281__vddio 500e-3
rj584 n128__vddio n282__vddio 500e-3
rj585 n124__vddio n283__vddio 500e-3
rj586 n120__vddio n284__vddio 500e-3
rj587 n116__vddio n285__vddio 500e-3
rj588 n112__vddio n286__vddio 500e-3
rj589 n108__vddio n287__vddio 500e-3
rj590 n104__vddio n288__vddio 500e-3
rj591 n100__vddio n289__vddio 500e-3
rj592 n96__vddio n290__vddio 500e-3
rj593 n92__vddio n291__vddio 500e-3
rj594 n88__vddio n292__vddio 500e-3
rj595 n84__vddio n293__vddio 500e-3
rj596 n80__vddio n294__vddio 500e-3
rj597 n76__vddio n295__vddio 500e-3
rj598 n72__vddio n296__vddio 500e-3
rj599 n68__vddio n297__vddio 500e-3
rj600 n64__vddio n298__vddio 500e-3
rj601 n60__vddio n299__vddio 500e-3
rj602 n56__vddio n300__vddio 500e-3
rj603 n52__vddio n301__vddio 500e-3
rj604 n396__vss n397__vss 414e-3
rj605 n397__vss n398__vss 327.1e-3
rj606 n398__vss n399__vss 334.4e-3
rj607 n399__vss n400__vss 327.1e-3
rj608 n400__vss n401__vss 327.1e-3
rj609 n401__vss n402__vss 334.4e-3
rj610 n402__vss n403__vss 327.1e-3
rj611 n403__vss n404__vss 327.1e-3
rj612 n404__vss n405__vss 334.4e-3
rj613 n405__vss n406__vss 327.1e-3
rj614 n406__vss n407__vss 327.1e-3
rj615 n407__vss n408__vss 327.1e-3
rj616 n408__vss n409__vss 327.1e-3
rj617 n409__vss n410__vss 327.1e-3
rj618 n410__vss n411__vss 334.4e-3
rj619 n411__vss n412__vss 327.1e-3
rj620 n412__vss n413__vss 327.1e-3
rj621 n413__vss n414__vss 334.4e-3
rj622 n414__vss n415__vss 327.1e-3
rj623 n415__vss n416__vss 327.1e-3
rj624 n416__vss n417__vss 334.4e-3
rj625 n417__vss n418__vss 327.1e-3
rj626 n418__vss n419__vss 327.1e-3
rj627 n419__vss n420__vss 341.6e-3
rj628 n420__vss n421__vss 327.1e-3
rj629 n421__vss n422__vss 334.4e-3
rj630 n422__vss n423__vss 327.1e-3
rj631 n423__vss n424__vss 327.1e-3
rj632 n424__vss n425__vss 334.4e-3
rj633 n425__vss n426__vss 327.1e-3
rj634 n426__vss n427__vss 327.1e-3
rj635 n427__vss n428__vss 334.4e-3
rj636 n428__vss n429__vss 327.1e-3
rj637 n429__vss n430__vss 327.1e-3
rj638 n430__vss n431__vss 327.1e-3
rj639 n431__vss n432__vss 327.1e-3
rj640 n432__vss n433__vss 327.1e-3
rj641 n433__vss n434__vss 334.4e-3
rj642 n434__vss n435__vss 327.1e-3
rj643 n435__vss n436__vss 327.1e-3
rj644 n436__vss n437__vss 339.2e-3
rj645 n437__vss n438__vss 327.1e-3
rj646 n438__vss n439__vss 327.1e-3
rj647 n439__vss n440__vss 334.4e-3
rj648 n440__vss n441__vss 327.1e-3
rj649 n441__vss n442__vss 327.1e-3
rj650 n442__vss n443__vss 332e-3
rj651 n443__vss n444__vss 334.4e-3
rj652 n444__vss n445__vss 327.1e-3
rj653 n445__vss n446__vss 327.8e-3
rj654 n446__vss n268__vss 3.7521
rj655 n395__vss n397__vss 500e-3
rj656 n393__vss n398__vss 500e-3
rj657 n391__vss n399__vss 500e-3
rj658 n389__vss n400__vss 500e-3
rj659 n387__vss n401__vss 500e-3
rj660 n385__vss n402__vss 500e-3
rj661 n383__vss n403__vss 500e-3
rj662 n381__vss n404__vss 500e-3
rj663 n379__vss n405__vss 500e-3
rj664 n377__vss n406__vss 500e-3
rj665 n375__vss n407__vss 500e-3
rj666 n373__vss n408__vss 500e-3
rj667 n371__vss n409__vss 500e-3
rj668 n369__vss n410__vss 500e-3
rj669 n367__vss n411__vss 500e-3
rj670 n365__vss n412__vss 500e-3
rj671 n363__vss n413__vss 500e-3
rj672 n361__vss n414__vss 500e-3
rj673 n359__vss n415__vss 500e-3
rj674 n357__vss n416__vss 500e-3
rj675 n355__vss n417__vss 500e-3
rj676 n353__vss n418__vss 500e-3
rj677 n351__vss n419__vss 500e-3
rj678 n349__vss n420__vss 500e-3
rj679 n347__vss n421__vss 500e-3
rj680 n345__vss n422__vss 500e-3
rj681 n343__vss n423__vss 500e-3
rj682 n341__vss n424__vss 500e-3
rj683 n338__vss n425__vss 500e-3
rj684 n336__vss n426__vss 500e-3
rj685 n334__vss n427__vss 500e-3
rj686 n332__vss n428__vss 500e-3
rj687 n330__vss n429__vss 500e-3
rj688 n328__vss n430__vss 500e-3
rj689 n326__vss n431__vss 500e-3
rj690 n324__vss n432__vss 500e-3
rj691 n322__vss n433__vss 500e-3
rj692 n320__vss n434__vss 500e-3
rj693 n318__vss n435__vss 500e-3
rj694 n316__vss n436__vss 500e-3
rj695 n314__vss n437__vss 500e-3
rj696 n312__vss n438__vss 500e-3
rj697 n310__vss n439__vss 500e-3
rj698 n308__vss n440__vss 500e-3
rj699 n306__vss n441__vss 500e-3
rj700 n304__vss n442__vss 500e-3
rj701 n302__vss n443__vss 500e-3
rj702 n300__vss n444__vss 500e-3
rj703 n298__vss n445__vss 500e-3
rj704 n296__vss n446__vss 500e-3
rk1 n5__i0__net2 n6__i0__net2 646.3e-3
rk2 n5__i0__net2 n7__i0__net2 75.4293
rk3 n4__i0__net2 n5__i0__net2 31
rk4 n11__clk n1__clk 503.3e-3
rk5 n8__i0__net1 n2__i0__net1 4.667e-3
rk6 n9__i0__net1 n10__i0__net1 4.667e-3
rk7 n8__i0__net1 n10__i0__net1 60.54e-3
rk9 n6__vdd n8__vdd 115.8e-3
rk10 n8__vdd n1__vdd 149.7e-3
rk11 n5__vdd n6__vdd 10.3333
rk12 n7__vdd n8__vdd 18.75
rk14 n6__vss n8__vss 117.6e-3
rk15 n8__vss n1__vss 199e-3
rk17 n5__vss n6__vss 25
rk18 n7__vss n8__vss 15.5
rk19 n5__clk n12__clk 1.1502
rk20 n8__i0__net2 i0__net2 3.292e-3
rk21 n9__i0__net2 n10__i0__net2 3.292e-3
rk22 n8__i0__net2 n10__i0__net2 17.03e-3
rk23 n4__clkb clkb 466.1e-3
rk25 n13__clk n8__clk 2.56e-3
rk26 n6__clkb n7__clkb 275.8e-3
rk27 n7__clkb n8__clkb 25.2482
rk28 n7__clkb n9__clkb 10.7078
rk29 n3__clk2 n9__clk2 165.7e-3
rk30 n9__clk2 n10__clk2 146e-3
rk31 n10__clk2 n11__clk2 31.1668
rk32 n9__clk2 n12__clk2 75.1143
rk33 n12__i0__net1 n13__i0__net1 75.126
rk34 n13__i0__net1 n15__i0__net1 287.7e-3
rk35 n15__i0__net1 n11__i0__net1 156.9e-3
rk36 n14__i0__net1 n15__i0__net1 31
rk37 n5__i0__net6 n6__i0__net6 650.3e-3
rk38 n5__i0__net6 n7__i0__net6 75.4569
rk39 n4__i0__net6 n5__i0__net6 31
rk40 n14__clk2 n5__clk2 503.3e-3
rk41 n8__i0__net4 n2__i0__net4 4.873e-3
rk42 n9__i0__net4 n10__i0__net4 4.873e-3
rk43 n8__i0__net4 n10__i0__net4 55.88e-3
rk44 n8__i0__net6 i0__net6 3.292e-3
rk45 n9__i0__net6 n10__i0__net6 3.292e-3
rk46 n8__i0__net6 n10__i0__net6 16.89e-3
rk47 n7__i0__net1 n16__i0__net1 458.6e-3
rk48 n16__i0__net1 n4__i0__net1 8.891e-3
rk49 n15__clk2 n8__clk2 2.56e-3
rk50 n3__i0__net3 n5__i0__net3 180.1e-3
rk51 n5__i0__net3 n6__i0__net3 75.1186
rk52 n5__i0__net3 n7__i0__net3 31.3216
rk53 n12__i0__net4 n13__i0__net4 75.1396
rk54 n13__i0__net4 n15__i0__net4 289.1e-3
rk55 n15__i0__net4 n11__i0__net4 151.9e-3
rk56 n13__i0__net4 n6__i0__net4 179.1e-3
rk57 n14__i0__net4 n15__i0__net4 31
rk58 n33__clk4 n34__clk4 31.1889
rk59 n34__clk4 n35__clk4 87.27e-3
rk60 n35__clk4 n36__clk4 75.1354
rk61 n35__clk4 n3__clk4 175.2e-3
rk62 n29__clk4b n31__clk4b 31.4057
rk63 n31__clk4b n32__clk4b 500e-3
rk64 n30__clk4b n31__clk4b 75
rk65 n5__i2__net1 n6__i2__net1 631.9e-3
rk66 n5__i2__net1 n7__i2__net1 75.4253
rk67 n4__i2__net1 n5__i2__net1 31
rk68 n5__i1__net1 n6__i1__net1 631.9e-3
rk69 n5__i1__net1 n7__i1__net1 75.426
rk70 n4__i1__net1 n5__i1__net1 31
rk71 n8__x2 n9__x2 2.477e-3
rk72 n2__x2 n9__x2 45
rk73 n14__vdd n15__vdd 16.1252
rk74 n8__x0 n9__x0 2.477e-3
rk75 n2__x0 n9__x0 45
rk76 n8__y2 n9__y2 3.259e-3
rk77 n2__y2 n8__y2 45
rk78 n41__clk4 n5__clk4 503.3e-3
rk79 n42__clk4 n7__clk4 503.3e-3
rk80 n16__vdd n17__vdd 16.1252
rk81 n7__vss n41__vss 20.7805
rk82 n41__vss vss 269.1e-3
rk83 vss n15__vss 182.8e-3
rk84 n41__vss n42__vss 460.3e-3
rk85 n42__vss n43__vss 37.5037
rk86 n4__yin0 yin0 4.867e-3
rk87 n2__yin0 n5__yin0 4.867e-3
rk88 n4__yin0 n5__yin0 50.57e-3
rk89 n4__xin0 xin0 6.489e-3
rk90 n2__xin0 n5__xin0 6.489e-3
rk91 n4__xin0 n5__xin0 43.35e-3
rk92 n8__y0 n9__y0 3.259e-3
rk93 n2__y0 n8__y0 45
rk94 n18__vdd n19__vdd 16.1174
rk95 n10__x2 n11__x2 3.375e-3
rk96 n6__x2 n12__x2 3.375e-3
rk97 n10__x2 n12__x2 11.72e-3
rk98 n8__i2__net1 i2__net1 6.489e-3
rk99 n8__i1__net1 i1__net1 6.489e-3
rk100 n6__clk4b n37__clk4b 290.2e-3
rk101 n37__clk4b clk4b 151e-3
rk102 n8__clk4b n38__clk4b 294.9e-3
rk103 n38__clk4b n3__clk4b 158.6e-3
rk104 n20__vdd n21__vdd 16.1174
rk105 n43__clk4 n10__clk4 2.56e-3
rk106 n44__clk4 n12__clk4 2.56e-3
rk107 n10__x0 n11__x0 3.375e-3
rk108 n6__x0 n12__x0 3.375e-3
rk109 n10__x0 n12__x0 11.72e-3
rk110 n10__y0 n12__y0 3.838e-3
rk111 n12__y0 n13__y0 75.4311
rk112 n11__y0 n12__y0 31
rk113 n13__x0 n15__x0 3.838e-3
rk114 n15__x0 n16__x0 75.4311
rk115 n14__x0 n15__x0 31
rk116 n2__i5__bbar n5__i5__bbar 662e-3
rk117 n5__i5__bbar n6__i5__bbar 38.1386
rk118 n4__i5__bbar n5__i5__bbar 15.5
rk119 n2__rst n17__rst 4.584e-3
rk120 n4__rst n18__rst 4.584e-3
rk121 n2__i3__bbar n5__i3__bbar 662e-3
rk122 n5__i3__bbar n6__i3__bbar 38.1386
rk123 n4__i3__bbar n5__i3__bbar 15.5
rk124 n2__i5__abar n5__i5__abar 1.4181
rk125 n5__i5__abar n6__i5__abar 38.123
rk126 n4__i5__abar n5__i5__abar 15.5
rk127 n2__i3__abar n5__i3__abar 1.4181
rk128 n5__i3__abar n6__i3__abar 38.123
rk129 n4__i3__abar n5__i3__abar 15.5
rk130 n44__vss n45__vss 38.0051
rk131 n10__y2 n11__y2 3.375e-3
rk132 n6__y2 n12__y2 3.375e-3
rk133 n10__y2 n12__y2 11.83e-3
rk134 n4__y1 n5__y1 75.6849
rk135 n8__x1 n9__x1 75.6849
rk136 n5__rst n19__rst 4.584e-3
rk137 n7__rst n20__rst 4.584e-3
rk138 n9__i2__net1 n10__i2__net1 31.6484
rk139 n9__i1__net1 n10__i1__net1 31.6484
rk140 n46__vss n47__vss 38.0051
rk141 n55__vdd n30__vdd 16.4949
rk142 n30__vdd n56__vdd 314.2e-3
rk143 n56__vdd n57__vdd 19.5099
rk144 n56__vdd n25__vdd 376.9e-3
rk145 i5__net3 n2__i5__net3 75.8394
rk146 n16__y0 n17__y0 3.375e-3
rk147 n6__y0 n18__y0 3.375e-3
rk148 n16__y0 n18__y0 11.83e-3
rk149 n58__vdd n31__vdd 16.4949
rk150 n31__vdd n59__vdd 224.9e-3
rk151 n59__vdd n60__vdd 19.6021
rk152 n59__vdd n26__vdd 42.58e-3
rk153 i3__net3 n2__i3__net3 75.8394
rk154 n2__i2__rstb n9__i2__rstb 122.3e-3
rk155 n9__i2__rstb n4__i2__rstb 5.631e-3
rk156 n2__i1__rstb n9__i1__rstb 122.3e-3
rk157 n9__i1__rstb n4__i1__rstb 5.631e-3
rk158 a2 n2__a2 15.7754
rk159 n2__a2 n3__a2 37.9585
rk160 n2__a2 n4__a2 962.5e-3
rk161 n5__i2__net3 n6__i2__net3 635.5e-3
rk162 n5__i2__net3 n7__i2__net3 75.4536
rk163 n4__i2__net3 n5__i2__net3 31
rk164 n5__i1__net3 n6__i1__net3 635.5e-3
rk165 n5__i1__net3 n7__i1__net3 75.4536
rk166 n4__i1__net3 n5__i1__net3 31
rk167 a0 n2__a0 15.7754
rk168 n2__a0 n3__a0 37.9585
rk169 n2__a0 n4__a0 950.7e-3
rk170 n45__clk4 n13__clk4 503.3e-3
rk171 n46__clk4 n15__clk4 503.3e-3
rk172 n4__yin1 yin1 6.489e-3
rk173 n2__yin1 n5__yin1 6.489e-3
rk174 n4__yin1 n5__yin1 61.4e-3
rk175 n4__xin1 xin1 4.867e-3
rk176 n2__xin1 n5__xin1 4.867e-3
rk177 n4__xin1 n5__xin1 46.69e-3
rk178 n8__i2__net3 i2__net3 6.489e-3
rk179 n8__i1__net3 i1__net3 6.489e-3
rk180 n14__clk4b n41__clk4b 281.7e-3
rk181 n41__clk4b n9__clk4b 147.7e-3
rk182 n16__clk4b n42__clk4b 281.7e-3
rk183 n42__clk4b n11__clk4b 147.7e-3
rk184 n47__clk4 n18__clk4 2.56e-3
rk185 n48__clk4 n20__clk4 2.56e-3
rk186 n13__y1 n14__y1 522.9e-3
rk187 n14__y1 n15__y1 31.2784
rk188 n14__y1 n17__y1 168e-3
rk189 n17__y1 n11__y1 59.07e-3
rk190 n16__y1 n17__y1 75
rk191 n13__x1 n14__x1 522.9e-3
rk192 n14__x1 n15__x1 31.2784
rk193 n14__x1 n17__x1 168e-3
rk194 n17__x1 n11__x1 59.07e-3
rk195 n16__x1 n17__x1 75
rk196 n5__i2__net4 n6__i2__net4 631.9e-3
rk197 n5__i2__net4 n7__i2__net4 75.4539
rk198 n4__i2__net4 n5__i2__net4 31
rk199 n5__i1__net4 n6__i1__net4 631.9e-3
rk200 n5__i1__net4 n7__i1__net4 75.4539
rk201 n4__i1__net4 n5__i1__net4 31
rk202 n49__clk4 n21__clk4 503.3e-3
rk203 n50__clk4 n23__clk4 503.3e-3
rk204 n4__yin2 yin2 4.867e-3
rk205 n2__yin2 n5__yin2 4.867e-3
rk206 n4__yin2 n5__yin2 61.4e-3
rk207 n4__xin2 xin2 5.678e-3
rk208 n2__xin2 n5__xin2 5.678e-3
rk209 n4__xin2 n5__xin2 36.86e-3
rk210 n8__i2__net4 n3__i2__net4 3.244e-3
rk211 n9__i2__net4 n10__i2__net4 3.244e-3
rk212 n8__i2__net4 n10__i2__net4 16.3e-3
rk213 n8__i1__net4 n3__i1__net4 3.244e-3
rk214 n9__i1__net4 n10__i1__net4 3.244e-3
rk215 n8__i1__net4 n10__i1__net4 16.3e-3
rk216 n22__clk4b n43__clk4b 285.1e-3
rk217 n43__clk4b n17__clk4b 147.7e-3
rk218 n8__x3 n9__x3 2.477e-3
rk219 n2__x3 n9__x3 45
rk220 n24__clk4b n44__clk4b 285.1e-3
rk221 n44__clk4b n19__clk4b 147.7e-3
rk222 n51__clk4 n52__clk4 1.392e-3
rk223 n26__clk4 n53__clk4 1.392e-3
rk224 n52__clk4 n53__clk4 10.24e-3
rk225 n54__clk4 n55__clk4 1.392e-3
rk226 n28__clk4 n56__clk4 1.392e-3
rk227 n55__clk4 n56__clk4 10.24e-3
rk228 n61__vdd n62__vdd 16.1252
rk229 n7__vss n68__vss 20.7684
rk230 n68__vss n69__vss 583.3e-3
rk231 n69__vss n70__vss 2.0268
rk232 n70__vss n7__vss 20.8063
rk233 n68__vss n71__vss 475.4e-3
rk234 n71__vss n72__vss 37.5025
rk235 n69__vss n50__vss 106.1e-3
rk236 n70__vss n48__vss 434.5e-3
rk237 n48__vss n73__vss 37.5037
rk238 n15__y2 n16__y2 75.2583
rk239 n16__y2 n17__y2 31.1458
rk240 n15__x2 n16__x2 75.2583
rk241 n16__x2 n17__x2 31.1458
rk242 n10__rst n29__rst 4.584e-3
rk243 n8__y3 n9__y3 3.259e-3
rk244 n2__y3 n8__y3 45
rk245 n12__rst n30__rst 4.584e-3
rk246 n10__i2__rstb n11__i2__rstb 3.132e-3
rk247 n6__i2__rstb n12__i2__rstb 3.132e-3
rk248 n10__i2__rstb n12__i2__rstb 18.42e-3
rk249 n10__i1__rstb n11__i1__rstb 3.132e-3
rk250 n6__i1__rstb n12__i1__rstb 3.132e-3
rk251 n10__i1__rstb n12__i1__rstb 18.42e-3
rk252 n63__vdd n64__vdd 16.1174
rk253 n5__i2__net2 n6__i2__net2 635.5e-3
rk254 n5__i2__net2 n7__i2__net2 75.4477
rk255 n4__i2__net2 n5__i2__net2 31
rk256 n10__x3 n11__x3 3.375e-3
rk257 n6__x3 n12__x3 3.375e-3
rk258 n10__x3 n12__x3 11.72e-3
rk259 n5__i1__net2 n6__i1__net2 635.5e-3
rk260 n5__i1__net2 n7__i1__net2 75.4477
rk261 n4__i1__net2 n5__i1__net2 31
rk262 n19__x1 n20__x1 2.477e-3
rk263 n2__x1 n20__x1 45
rk264 n70__vdd n71__vdd 16.1252
rk265 n7__vss n74__vss 20.7805
rk266 n74__vss n51__vss 1.0706
rk267 n74__vss n75__vss 453e-3
rk268 n75__vss n76__vss 37.5037
rk269 n57__clk4 n29__clk4 503.3e-3
rk270 n58__clk4 n31__clk4 503.3e-3
rk271 n2__i6__bbar n5__i6__bbar 662e-3
rk272 n5__i6__bbar n6__i6__bbar 38.1393
rk273 n4__i6__bbar n5__i6__bbar 15.5
rk274 n4__yin3 yin3 4.867e-3
rk275 n2__yin3 n5__yin3 4.867e-3
rk276 n4__yin3 n5__yin3 17.2e-3
rk277 n4__xin3 xin3 5.678e-3
rk278 n2__xin3 n5__xin3 5.678e-3
rk279 n4__xin3 n5__xin3 19.66e-3
rk280 n19__y1 n20__y1 3.259e-3
rk281 n2__y1 n19__y1 45
rk282 n2__i6__abar n5__i6__abar 1.4181
rk283 n5__i6__abar n6__i6__abar 38.123
rk284 n4__i6__abar n5__i6__abar 15.5
rk285 n77__vss n78__vss 38.0051
rk286 n10__y3 n11__y3 3.375e-3
rk287 n6__y3 n12__y3 3.375e-3
rk288 n10__y3 n12__y3 11.83e-3
rk289 n8__i2__net2 i2__net2 6.489e-3
rk290 n72__vdd n73__vdd 16.1174
rk291 n8__i1__net2 i1__net2 6.489e-3
rk292 n34__clk4b n45__clk4b 281.7e-3
rk293 n45__clk4b n25__clk4b 147.7e-3
rk294 n36__clk4b n46__clk4b 281.7e-3
rk295 n46__clk4b n27__clk4b 147.7e-3
rk296 n59__clk4 n38__clk4 2.56e-3
rk297 n21__x1 n22__x1 3.375e-3
rk298 n6__x1 n23__x1 3.375e-3
rk299 n21__x1 n23__x1 11.72e-3
rk300 n60__clk4 n40__clk4 2.56e-3
rk301 n74__vdd n75__vdd 16.3364
rk302 n75__vdd n65__vdd 173e-3
rk303 n65__vdd n76__vdd 19.8131
rk304 n75__vdd n68__vdd 124.9e-3
rk305 i6__net3 n2__i6__net3 75.8088
rk306 n2__i4__bbar n5__i4__bbar 662e-3
rk307 n5__i4__bbar n6__i4__bbar 38.1386
rk308 n4__i4__bbar n5__i4__bbar 15.5
rk309 n16__y3 n14__y3 75.1404
rk310 n14__y3 n18__y3 4.657e-3
rk311 n14__y3 n19__y3 31.4301
rk312 n17__y3 n18__y3 75
rk313 n13__i2__net4 n11__i2__net4 31.1484
rk314 n16__x3 n15__x3 75.1404
rk315 n15__x3 n18__x3 4.657e-3
rk316 n15__x3 n19__x3 31.4301
rk317 n17__x3 n18__x3 75
rk318 n13__i1__net4 n11__i1__net4 31.1484
rk319 n2__i4__abar n5__i4__abar 1.4181
rk320 n5__i4__abar n6__i4__abar 38.123
rk321 n4__i4__abar n5__i4__abar 15.5
rk322 n96__vdd n97__vdd 31.8842
rk323 n97__vdd n98__vdd 447e-3
rk324 n98__vdd n99__vdd 472.7e-3
rk325 n99__vdd n100__vdd 769.8e-3
rk326 n100__vdd n101__vdd 447e-3
rk327 n101__vdd n102__vdd 323.1e-3
rk328 n102__vdd n103__vdd 462.9e-3
rk329 n103__vdd n29__vdd 47.52e-3
rk330 n97__vdd n104__vdd 31.278
rk331 n98__vdd n105__vdd 31.262
rk332 n99__vdd n106__vdd 31.2787
rk333 n100__vdd n107__vdd 31.278
rk334 n101__vdd n108__vdd 31.2861
rk335 n102__vdd n109__vdd 25.2409
rk336 n103__vdd n110__vdd 31.2887
rk337 n79__vss n80__vss 75.7757
rk338 n80__vss n81__vss 443.5e-3
rk339 n81__vss n82__vss 440.3e-3
rk340 n82__vss n83__vss 711.8e-3
rk341 n83__vss n84__vss 445.6e-3
rk342 n84__vss n85__vss 347.7e-3
rk343 n85__vss n86__vss 440.3e-3
rk344 n86__vss n20__vss 843.3e-3
rk345 n80__vss n87__vss 75.2014
rk346 n81__vss n88__vss 75.2033
rk347 n82__vss n89__vss 75.2014
rk348 n83__vss n90__vss 75.2014
rk349 n84__vss n7__vss 20.85
rk350 n85__vss n91__vss 75.2212
rk351 n86__vss n92__vss 75.2014
rk352 n111__vdd n112__vdd 31.8842
rk353 n112__vdd n113__vdd 213.7e-3
rk354 n113__vdd n114__vdd 274.1e-3
rk355 n114__vdd n115__vdd 472.7e-3
rk356 n115__vdd n116__vdd 769.8e-3
rk357 n116__vdd n117__vdd 447e-3
rk358 n117__vdd n118__vdd 323.1e-3
rk359 n118__vdd n22__vdd 482.4e-3
rk360 n112__vdd n119__vdd 31.278
rk361 n113__vdd n66__vdd 61.2e-3
rk362 n114__vdd n120__vdd 31.262
rk363 n115__vdd n121__vdd 31.2787
rk364 n116__vdd n122__vdd 31.278
rk365 n117__vdd n123__vdd 31.2861
rk366 n118__vdd n124__vdd 25.2409
rk367 n22__vdd n125__vdd 31.2895
rk368 n22__vdd n126__vdd 916e-3
rk369 n126__vdd n127__vdd 79.83e-3
rk370 n127__vdd n128__vdd 31.1607
rk371 n126__vdd n129__vdd 308.7e-3
rk372 n129__vdd n130__vdd 31.2565
rk373 n127__vdd n131__vdd 31.4702
rk374 n129__vdd n132__vdd 546.2e-3
rk375 n132__vdd n133__vdd 31.3511
rk376 n132__vdd n134__vdd 519.1e-3
rk377 n134__vdd n124__vdd 25.2371
rk378 n134__vdd n135__vdd 303.6e-3
rk379 n135__vdd n136__vdd 31.2622
rk380 n135__vdd n137__vdd 31.7532
rk381 n93__vss n94__vss 75.7757
rk382 n94__vss n95__vss 443.5e-3
rk383 n95__vss n96__vss 440.3e-3
rk384 n96__vss n97__vss 711.8e-3
rk385 n97__vss n98__vss 445.6e-3
rk386 n98__vss n99__vss 347.7e-3
rk387 n99__vss n100__vss 442.8e-3
rk388 n100__vss n17__vss 895.4e-3
rk389 n17__vss n101__vss 94.88e-3
rk390 n101__vss n102__vss 314.8e-3
rk391 n102__vss n103__vss 470.5e-3
rk392 n103__vss n104__vss 479.7e-3
rk393 n104__vss n105__vss 329.9e-3
rk394 n105__vss n106__vss 75.5773
rk395 n94__vss n107__vss 75.2014
rk396 n95__vss n108__vss 75.2033
rk397 n96__vss n109__vss 75.2014
rk398 n97__vss n110__vss 75.2014
rk399 n98__vss n7__vss 20.85
rk400 n99__vss n111__vss 75.2212
rk401 n100__vss n112__vss 75.2014
rk402 n101__vss n113__vss 75.1101
rk403 n101__vss n114__vss 75.4509
rk404 n102__vss n115__vss 75.0896
rk405 n103__vss n116__vss 75.0963
rk406 n104__vss n7__vss 20.7341
rk407 n105__vss n117__vss 75.0911
rk408 n118__vss n119__vss 38.0051
rk409 n23__rst n36__rst 137.9e-3
rk410 n36__rst n14__rst 2.815e-3
rk411 n27__rst n43__rst 137.9e-3
rk412 n43__rst n16__rst 2.815e-3
rk413 n22__y1 n23__y1 3.375e-3
rk414 n9__y1 n24__y1 3.375e-3
rk415 n22__y1 n24__y1 11.83e-3
rk416 n13__i2__rstb n14__i2__rstb 31.1643
rk417 n14__i2__rstb n7__i2__rstb 149.1e-3
rk418 n7__i2__rstb n15__i2__rstb 508.4e-3
rk419 n14__i2__rstb n16__i2__rstb 75.2695
rk420 n13__i1__rstb n14__i1__rstb 31.1643
rk421 n14__i1__rstb n7__i1__rstb 149.1e-3
rk422 n7__i1__rstb n15__i1__rstb 508.4e-3
rk423 n14__i1__rstb n16__i1__rstb 75.2695
rk424 n138__vdd n79__vdd 16.4712
rk425 n79__vdd n78__vdd 366.2e-3
rk426 n78__vdd n139__vdd 19.3881
rk427 i4__net3 n2__i4__net3 75.8199
rk428 n9__a1 n10__a1 15.7754
rk429 n10__a1 n11__a1 37.9585
rk430 n10__a1 n12__a1 956.2e-3
rk431 n9__a3 n10__a3 1.7453
rk432 n10__a3 n11__a3 37.9592
rk433 n10__a3 n12__a3 15.7754
rk434 n13__a2 n14__a2 2.399e-3
rk435 n6__a2 n14__a2 45
rk436 n13__a0 n14__a0 2.399e-3
rk437 n6__a0 n14__a0 45
rk438 n4__i8__net51 n5__i8__net51 75.5
rk439 n4__i7__net51 n5__i7__net51 75.5
rk440 n13__a3 n2__a3 45.5072
rk441 n13__a1 n2__a1 45.5072
rk442 i8__net49 n2__i8__net49 31.7999
rk444 n7__i8__net51 n8__i8__net51 15.5818
rk445 n7__i8__net51 n9__i8__net51 177.5e-3
rk446 n9__i8__net51 n2__i8__net51 45.0028
rk447 i7__net49 n2__i7__net49 31.7999
rk449 n7__i7__net51 n8__i7__net51 15.5818
rk450 n7__i7__net51 n9__i7__net51 177.5e-3
rk451 n9__i7__net51 n2__i7__net51 45.0028
rk452 n9__s1 n10__s1 16.1074
rk453 n10__s1 n11__s1 411.7e-3
rk454 n11__s1 n12__s1 38.163
rk455 n11__s1 n13__s1 75.1591
rk456 n9__s0 n10__s0 16.0015
rk457 n10__s0 n11__s0 522e-3
rk458 n11__s0 n12__s0 38.163
rk459 n11__s0 n13__s0 75.1591
rk460 n17__c1 n18__c1 31.9138
rk461 n18__c1 n19__c1 75.187
rk462 n18__c0 n19__c0 542.2e-3
rk463 n18__c0 n20__c0 76.119
rk464 n17__c0 n18__c0 31
rk465 n15__a2 n16__a2 4.224e-3
rk466 n11__a2 n15__a2 45
rk467 n15__a0 n16__a0 4.224e-3
rk468 n11__a0 n15__a0 45
rk469 n4__i8__carry_bar n5__i8__carry_bar 31.5867
rk470 n5__i8__carry_bar n2__i8__carry_bar 45.2091
rk471 n5__i8__carry_bar n6__i8__carry_bar 38.2157
rk472 n4__i7__carry_bar n5__i7__carry_bar 31.5867
rk473 n5__i7__carry_bar n2__i7__carry_bar 45.2091
rk474 n5__i7__carry_bar n6__i7__carry_bar 38.2157
rk475 n139__vss n140__vss 38.417
rk476 n140__vss n141__vss 314e-3
rk477 n141__vss n142__vss 314e-3
rk478 n142__vss n143__vss 288.7e-3
rk479 n143__vss n144__vss 273e-3
rk480 n144__vss n121__vss 300.3e-3
rk481 n140__vss n145__vss 75.4558
rk482 n141__vss n146__vss 75.4558
rk483 n142__vss n148__vss 149.6e-3
rk484 n148__vss n149__vss 37.7817
rk485 n143__vss n150__vss 75.1496
rk486 n144__vss n7__vss 20.9794
rk487 n147__vss n148__vss 75
rk488 n152__vdd n153__vdd 31.529
rk489 n153__vdd n154__vdd 184.6e-3
rk490 n154__vdd n155__vdd 528e-3
rk491 n155__vdd n156__vdd 338.5e-3
rk492 n156__vdd n157__vdd 896.1e-3
rk493 n157__vdd n158__vdd 518.3e-3
rk494 n158__vdd n160__vdd 171.2e-3
rk495 n153__vdd n161__vdd 31.2485
rk496 n154__vdd n162__vdd 31.2485
rk497 n155__vdd n151__vdd 33.55e-3
rk498 n156__vdd n163__vdd 15.833
rk499 n157__vdd n164__vdd 15.775
rk500 n158__vdd n165__vdd 25.1851
rk502 n159__vdd n160__vdd 15.5
rk503 n15__a3 n16__a3 11.77e-3
rk504 n7__a3 n15__a3 45
rk505 n14__a3 n16__a3 500e-3
rk506 n167__vdd n168__vdd 31.529
rk507 n168__vdd n169__vdd 184.6e-3
rk508 n169__vdd n170__vdd 522.4e-3
rk509 n170__vdd n171__vdd 105.7e-3
rk510 n171__vdd n172__vdd 896.1e-3
rk511 n172__vdd n173__vdd 518.3e-3
rk512 n173__vdd n175__vdd 171.2e-3
rk513 n168__vdd n176__vdd 31.2485
rk514 n169__vdd n177__vdd 31.2499
rk515 n170__vdd n148__vdd 220.1e-3
rk516 n171__vdd n178__vdd 15.8327
rk517 n172__vdd n179__vdd 15.775
rk518 n173__vdd n180__vdd 25.1851
rk520 n174__vdd n175__vdd 15.5
rk521 n14__a1 n15__a1 11.77e-3
rk522 n7__a1 n14__a1 45
rk523 n14__s0 n15__s0 2.399e-3
rk524 n2__s0 n15__s0 45
rk525 n12__i10__net116 n9__i10__net116 11.86e-3
rk526 n9__i10__net116 n13__i10__net116 15.5211
rk527 n11__i10__net116 n12__i10__net116 7.75
rk528 n4__i9__net51 n5__i9__net51 75.5
rk529 n16__s1 n2__s1 45.5072
rk531 n2__i10__net124 n4__i10__net124 5.631e-3
rk533 n3__i10__net124 n4__i10__net124 18.75
rk535 n2__i10__net115 n4__i10__net115 45.05e-3
rk536 n3__i10__net115 n4__i10__net115 7.75
rk537 i9__net49 n2__i9__net49 31.7999
rk539 n7__i9__net51 n8__i9__net51 15.5818
rk540 n7__i9__net51 n9__i9__net51 177.5e-3
rk541 n9__i9__net51 n2__i9__net51 45.0028
rk543 i10__net115 n8__i10__net115 45.05e-3
rk544 n7__i10__net115 n8__i10__net115 7.75
rk546 i10__net124 n9__i10__net124 5.631e-3
rk548 n8__i10__net124 n9__i10__net124 18.75
rk549 r0 n2__r0 16.2255
rk550 n2__r0 n3__r0 281.1e-3
rk551 n3__r0 n4__r0 38.163
rk552 n3__r0 n5__r0 75.1591
rk553 n7__i10__net114 n8__i10__net114 16.3867
rk554 n9__i10__net114 n10__i10__net114 38.2097
rk555 n15__i10__net116 n16__i10__net116 31.66e-3
rk556 n16__i10__net116 n17__i10__net116 37.5317
rk557 n16__i10__net116 n10__i10__net116 102.2e-3
rk558 n10__i10__net116 n18__i10__net116 696.5e-3
rk559 n18__i10__net116 n3__i10__net116 25.61e-3
rk560 n14__i10__net116 n15__i10__net116 18.75
rk561 n14__net12 n15__net12 542.2e-3
rk562 n14__net12 n16__net12 76.1062
rk563 n13__net12 n14__net12 31
rk565 n3__i10__net122 n4__i10__net122 5.631e-3
rk567 n2__i10__net122 n3__i10__net122 15.5
rk568 i10__net125 n3__i10__net125 10.61e-3
rk569 n2__i10__net125 n3__i10__net125 37.5
rk570 n16__s0 n17__s0 4.224e-3
rk571 n7__s0 n16__s0 45
rk572 n4__i10__net125 n6__i10__net125 10.61e-3
rk573 n5__i10__net125 n6__i10__net125 37.5
rk575 n8__i10__net122 i10__net122 5.631e-3
rk577 n7__i10__net122 n8__i10__net122 15.5
rk578 n4__i9__carry_bar n5__i9__carry_bar 31.5867
rk579 n5__i9__carry_bar n2__i9__carry_bar 45.2091
rk580 n5__i9__carry_bar n6__i9__carry_bar 38.2157
rk581 n191__vdd n192__vdd 31.4249
rk582 n192__vdd n193__vdd 124.6e-3
rk583 n193__vdd n194__vdd 184.6e-3
rk584 n194__vdd n195__vdd 607.6e-3
rk585 n195__vdd n196__vdd 896.1e-3
rk586 n196__vdd n197__vdd 518.3e-3
rk587 n197__vdd n199__vdd 171.2e-3
rk588 n192__vdd n187__vdd 221.9e-3
rk589 n193__vdd n200__vdd 31.2485
rk590 n194__vdd n201__vdd 31.2499
rk591 n195__vdd n202__vdd 15.8327
rk592 n196__vdd n203__vdd 15.775
rk593 n197__vdd n180__vdd 25.1851
rk595 n198__vdd n199__vdd 15.5
rk596 n17__s1 n18__s1 11.77e-3
rk597 n7__s1 n17__s1 45
rk598 n169__vss n170__vss 38.3521
rk599 n170__vss n171__vss 300.6e-3
rk600 n171__vss n172__vss 293.4e-3
rk601 n172__vss n158__vss 59.12e-3
rk602 n158__vss n173__vss 193.1e-3
rk603 n173__vss n174__vss 261.5e-3
rk604 n174__vss n175__vss 287.3e-3
rk605 n175__vss n176__vss 437.7e-3
rk606 n176__vss n177__vss 314e-3
rk607 n177__vss n178__vss 314e-3
rk608 n178__vss n179__vss 288.7e-3
rk609 n179__vss n180__vss 273e-3
rk610 n180__vss n122__vss 369.8e-3
rk611 n170__vss n181__vss 75.4546
rk612 n171__vss n182__vss 75.4546
rk613 n172__vss n184__vss 149.9e-3
rk614 n184__vss n185__vss 37.7817
rk615 n173__vss n186__vss 75.1487
rk616 n174__vss n7__vss 20.9774
rk617 n175__vss n187__vss 37.9183
rk618 n176__vss n188__vss 75.4558
rk619 n177__vss n189__vss 75.4558
rk620 n178__vss n191__vss 149.6e-3
rk621 n191__vss n192__vss 37.7817
rk622 n179__vss n193__vss 75.1496
rk623 n180__vss n7__vss 20.9794
rk624 n183__vss n184__vss 75
rk625 n190__vss n191__vss 75
rk626 n11__i10__net114 n12__i10__net114 10.9893
rk627 n13__i10__net114 n14__i10__net114 25.6679
rk628 n11__net12 n7__net12 569.9e-3
rk629 n7__net12 n3__net12 745.8e-3
rk630 n3__net12 n17__net12 551.8e-3
rk631 n15__c1 n11__c1 697.8e-3
rk632 n11__c1 n7__c1 728.4e-3
rk633 n7__c1 n3__c1 714.5e-3
rk634 n3__c1 n20__c1 289.4e-3
rk635 n15__c0 n11__c0 605.4e-3
rk636 n11__c0 n7__c0 921.9e-3
rk637 n7__c0 n3__c0 622.3e-3
rk638 n3__c0 n21__c0 2.3102
rk639 i10__net114 n16__i10__net114 184.9e-3
rk640 n6__i10__net114 n17__i10__net114 126.1e-3
rk641 r1 n2__r1 31.3488
rk642 n2__r1 n3__r1 75.299
rk643 n19__i10__net116 n7__i10__net116 3.375e-3
rk645 n208__vdd n209__vdd 800.3e-3
rk646 n209__vdd n210__vdd 317.2e-3
rk647 n210__vdd n211__vdd 175.1e-3
rk648 n211__vdd n212__vdd 664.2e-3
rk649 n212__vdd n213__vdd 244.3e-3
rk650 n213__vdd n214__vdd 580.3e-3
rk651 n214__vdd n215__vdd 704.4e-3
rk653 n209__vdd n217__vdd 31.6375
rk654 n210__vdd n218__vdd 31.6774
rk655 n211__vdd n219__vdd 10.8435
rk656 n212__vdd n220__vdd 16.0787
rk657 n212__vdd n186__vdd 52.27e-3
rk658 n213__vdd n221__vdd 16.0905
rk659 n214__vdd n222__vdd 8.2269
rk660 n215__vdd n223__vdd 16.0568
rk661 n165__vdd n208__vdd 12.5
rk662 n194__vss n195__vss 75.3359
rk663 n195__vss n196__vss 325.7e-3
rk664 n196__vss n197__vss 175.1e-3
rk665 n197__vss n198__vss 578.5e-3
rk666 n198__vss n199__vss 279.3e-3
rk667 n199__vss n200__vss 590.5e-3
rk668 n200__vss n157__vss 197.1e-3
rk669 n157__vss n201__vss 491.2e-3
rk671 n195__vss n7__vss 12.9394
rk672 n196__vss n203__vss 75.3642
rk673 n197__vss n204__vss 25.2728
rk674 n198__vss n205__vss 37.8022
rk675 n199__vss n206__vss 37.8127
rk676 n200__vss n207__vss 18.9418
rk677 n201__vss n208__vss 37.7832
rk678 n4__r1 n5__r1 1.0762
rk679 r2 n2__r2 596.5e-3
rk680 n2__r2 n3__r2 75.1637
rk681 n2__r2 n4__r2 31.5079
rk682 n72__clk4 n73__clk4 1.688e-3
rk683 n70__clk4 n73__clk4 45
rk684 n5__i14__i7__net1 n6__i14__i7__net1 75.5017
rk685 n20__clk2 n21__clk2 1.765e-3
rk686 n18__clk2 n21__clk2 45
rk687 n7__i14__i7__net1 n8__i14__i7__net1 16.1187
rk688 n2__i14__i3__rstb n3__i14__i3__rstb 156.6e-3
rk689 n3__i14__i3__rstb n4__i14__i3__rstb 75.2698
rk690 n3__i14__i3__rstb n5__i14__i3__rstb 31.1638
rk691 n3__i14__i7__net1 n9__i14__i7__net1 500e-3
rk692 n49__rst n63__rst 142.2e-3
rk693 n63__rst n45__rst 2.329e-3
rk694 n25__i14__shift n26__i14__shift 528.5e-3
rk695 n26__i14__shift n27__i14__shift 75.2374
rk696 n26__i14__shift n28__i14__shift 31.2111
rk697 i14__net9 n2__i14__net9 31.1969
rk698 n2__i14__net9 n4__i14__net9 215.8e-3
rk699 n4__i14__net9 n5__i14__net9 75.1653
rk700 n3__i14__net9 n4__i14__net9 75
rk701 n15__clk n27__clk 2.56e-3
rk702 n4__i14__i3__net5 n5__i14__i3__net5 31.5125
rk703 n5__i14__i3__net5 n2__i14__i3__net5 3.128e-3
rk704 n228__vdd n230__vdd 31.2409
rk705 n230__vdd n231__vdd 436e-3
rk706 n231__vdd n232__vdd 130.8e-3
rk707 n232__vdd n233__vdd 31.2666
rk708 n229__vdd n230__vdd 25
rk709 n29__clk n18__clk 503.3e-3
rk710 n15__clkb n24__clkb 164.8e-3
rk711 n24__clkb n12__clkb 275.1e-3
rk712 n7__i14__i3__net5 n8__i14__i3__net5 75.4253
rk713 n7__i14__i3__net5 n9__i14__i3__net5 631.9e-3
rk714 n6__i14__i3__net5 n7__i14__i3__net5 31
rk715 n3__i14__shift n29__i14__shift 502.5e-3
rk716 n217__vss n218__vss 75.4027
rk717 n218__vss n219__vss 31.0851
rk718 n2__i14__i4__rstb n3__i14__i4__rstb 157e-3
rk719 n3__i14__i4__rstb n4__i14__i4__rstb 75.2698
rk720 n3__i14__i4__rstb n5__i14__i4__rstb 31.1638
rk721 n2__i14__i0__net1 n5__i14__i0__net1 503.4e-3
rk722 n6__i14__shift n30__i14__shift 3.371e-3
rk723 n55__rst n51__rst 146.1e-3
rk725 n8__i14__net2 n6__i14__net2 31.1605
rk726 n6__i14__net2 n9__i14__net2 75.3236
rk727 i14__net2 n7__i14__net2 854.4e-3
rk728 n4__i14__i0__net1 n8__i14__i0__net1 453.1e-3
rk729 n8__i14__i0__net1 n6__i14__i0__net1 261e-3
rk730 n6__i14__i0__net1 n9__i14__i0__net1 31.1737
rk731 n7__i14__i0__net1 n8__i14__i0__net1 75
rk732 n31__i14__shift n7__i14__shift 2.832e-3
rk733 i14__net15 n2__i14__net15 31.1969
rk734 n2__i14__net15 n4__i14__net15 215.8e-3
rk735 n4__i14__net15 n5__i14__net15 75.1653
rk736 n3__i14__net15 n4__i14__net15 75
rk737 n6__r2 n7__r2 31.1364
rk738 n7__r2 n8__r2 75.4102
rk739 n19__clk n35__clk 2.56e-3
rk740 n4__i14__i4__net5 n5__i14__i4__net5 31.5125
rk741 n5__i14__i4__net5 n2__i14__i4__net5 3.128e-3
rk742 n32__i14__shift n11__i14__shift 502e-3
rk743 n249__vdd n250__vdd 31.2524
rk744 n250__vdd n248__vdd 59.98e-3
rk745 n250__vdd n251__vdd 586.5e-3
rk746 n251__vdd n252__vdd 31.2666
rk747 n229__vdd n250__vdd 25
rk748 n36__clk n22__clk 503.3e-3
rk749 n19__clkb n25__clkb 164.8e-3
rk750 n25__clkb n16__clkb 275.1e-3
rk751 n7__i14__net9 n8__i14__net9 31.1786
rk752 n8__i14__net9 n9__i14__net9 75.3399
rk753 n4__i14__net8 i14__net8 772e-3
rk754 n14__i14__shift n33__i14__shift 3.371e-3
rk755 n2__i14__i1__net1 n5__i14__i1__net1 503.4e-3
rk756 n7__i14__i4__net5 n8__i14__i4__net5 75.4253
rk757 n7__i14__i4__net5 n9__i14__i4__net5 631.9e-3
rk758 n6__i14__i4__net5 n7__i14__i4__net5 31
rk759 n5__i14__net8 n6__i14__net8 31.1619
rk760 n6__i14__net8 n7__i14__net8 75.3242
rk761 n4__i14__i1__net1 n7__i14__i1__net1 458e-3
rk762 n7__i14__i1__net1 n8__i14__i1__net1 273.6e-3
rk763 n8__i14__i1__net1 n9__i14__i1__net1 31.1837
rk764 n6__i14__i1__net1 n7__i14__i1__net1 75
rk765 n34__i14__shift n15__i14__shift 2.832e-3
rk766 n8__r1 n9__r1 31.1364
rk767 n9__r1 n10__r1 75.4102
rk768 n2__i14__i5__rstb n3__i14__i5__rstb 156.6e-3
rk769 n3__i14__i5__rstb n4__i14__i5__rstb 75.2698
rk770 n3__i14__i5__rstb n5__i14__i5__rstb 31.1638
rk771 n253__vdd n255__vdd 31.4212
rk772 n255__vdd n256__vdd 615.3e-3
rk773 n256__vdd n257__vdd 760.5e-3
rk774 n256__vdd n258__vdd 31.2738
rk775 n257__vdd n259__vdd 31.302
rk776 n257__vdd n260__vdd 455.7e-3
rk777 n260__vdd n236__vdd 53.9e-3
rk778 n260__vdd n262__vdd 249.5e-3
rk779 n262__vdd n263__vdd 31.2688
rk780 n260__vdd n234__vdd 829e-3
rk781 n262__vdd n264__vdd 16.2454
rk782 n254__vdd n255__vdd 18.75
rk783 n254__vdd n257__vdd 9.375
rk784 n261__vdd n262__vdd 12.5
rk785 n35__i14__shift n19__i14__shift 502e-3
rk786 n61__rst n70__rst 142.2e-3
rk787 n70__rst n57__rst 2.329e-3
rk788 n6__serial_out n7__serial_out 31.2685
rk789 n7__serial_out n9__serial_out 136.7e-3
rk790 n9__serial_out n10__serial_out 75.1667
rk791 n8__serial_out n9__serial_out 75
rk792 n7__i14__net15 n8__i14__net15 31.1786
rk793 n8__i14__net15 n9__i14__net15 75.3399
rk794 n22__i14__shift n36__i14__shift 3.371e-3
rk795 n2__i14__i2__net1 n5__i14__i2__net1 503.4e-3
rk796 n23__clk n38__clk 2.56e-3
rk797 n4__i14__i5__net5 n5__i14__i5__net5 31.5125
rk798 n5__i14__i5__net5 n2__i14__i5__net5 3.128e-3
rk799 n4__i14__net14 n5__i14__net14 31.1618
rk800 n5__i14__net14 n6__i14__net14 75.3235
rk801 n223__vss n224__vss 75.5066
rk802 n224__vss n225__vss 199.3e-3
rk803 n225__vss n226__vss 587.4e-3
rk804 n226__vss n227__vss 339.3e-3
rk805 n227__vss n228__vss 199.3e-3
rk806 n228__vss n229__vss 587.4e-3
rk807 n229__vss n230__vss 339.3e-3
rk808 n230__vss n231__vss 199.3e-3
rk809 n231__vss n209__vss 378.2e-3
rk811 n225__vss n233__vss 75.1633
rk812 n226__vss n234__vss 75.1635
rk813 n228__vss n235__vss 75.1633
rk814 n229__vss n236__vss 75.1635
rk815 n231__vss n237__vss 75.1633
rk816 n209__vss n238__vss 689.3e-3
rk817 n238__vss n239__vss 622.7e-3
rk818 n239__vss n240__vss 75.2175
rk819 n239__vss n241__vss 253.5e-3
rk820 n241__vss n242__vss 75.1987
rk821 n241__vss n243__vss 172e-3
rk822 n243__vss n244__vss 75.1976
rk823 n243__vss n245__vss 673.9e-3
rk824 n245__vss n246__vss 75.4569
rk825 n245__vss n221__vss 422.5e-3
rk826 n221__vss n247__vss 476.2e-3
rk827 n247__vss n248__vss 75.2945
rk828 n247__vss n249__vss 76.0373
rk829 n7__vss n224__vss 20.6667
rk830 n7__vss n227__vss 20.6667
rk831 n7__vss n230__vss 20.6667
rk832 n7__vss n238__vss 4.1333
rk833 n266__vdd n267__vdd 31.2524
rk834 n267__vdd n265__vdd 57.58e-3
rk835 n267__vdd n268__vdd 31.8853
rk836 n229__vdd n267__vdd 25
rk837 n4__i14__i2__net1 n8__i14__i2__net1 458e-3
rk838 n8__i14__i2__net1 n6__i14__i2__net1 273.6e-3
rk839 n6__i14__i2__net1 n9__i14__i2__net1 31.1837
rk840 n7__i14__i2__net1 n8__i14__i2__net1 75
rk841 n37__i14__shift n23__i14__shift 2.832e-3
rk842 n10__r0 n12__r0 75.5357
rk843 n12__r0 n13__r0 578e-3
rk844 n11__r0 n12__r0 31
rk845 i14__net14 n8__i14__net14 306.8e-3
rk846 n39__clk n26__clk 503.3e-3
rk847 n23__clkb n26__clkb 164.8e-3
rk848 n26__clkb n20__clkb 275.1e-3
rk849 n7__i14__i5__net5 n8__i14__i5__net5 75.4253
rk850 n7__i14__i5__net5 n9__i14__i5__net5 631.9e-3
rk851 n6__i14__i5__net5 n7__i14__i5__net5 31
rk853 n3__vddio n5__vddio 542.4e-3
rk854 n5__vddio n6__vddio 252.3e-3
rk855 n2__vddio n3__vddio 12.4
rk856 n4__vddio n5__vddio 25
rk857 n4__i11__net1 n5__i11__net1 531e-3
rk858 n4__i11__net1 n6__i11__net1 75.3087
rk859 n3__i11__net1 n4__i11__net1 31
rk860 net5 n3__net5 334.4e-3
rk861 n3__net5 n4__net5 4.9931
rk862 n3__net5 n5__net5 12.8501
rk863 n4__serial_out n12__serial_out 216.8e-3
rk864 n12__serial_out serial_out 42.02e-3
rk865 n7__i11__net1 i11__net1 2.512e-3
rk867 n273__vdd n270__vdd 65.2e-3
rk868 n270__vdd n275__vdd 58.21e-3
rk870 n272__vdd n273__vdd 25
rk871 n274__vdd n275__vdd 31
rk872 n7__vss n250__vss 20.7855
rk873 n250__vss n253__vss 58.21e-3
rk874 n253__vss n254__vss 6.311
rk875 n252__vss n253__vss 75
rk876 n6__r_in n7__r_in 12.7606
rk877 n7__r_in r_in 334.4e-3
rk878 n7__r_in n8__r_in 229.8e-3
rk879 n8__r_in n9__r_in 4.8731
rk880 n8__r_in n3__r_in 47.1462
rk881 n31__i12__net2 n32__i12__net2 8.8107
rk882 n32__i12__net2 n33__i12__net2 1.5153
rk883 n33__i12__net2 n34__i12__net2 518.3e-3
rk885 n31__i12__net2 n32__i12__net2 3.1
rk886 n31__i12__net2 n33__i12__net2 3.1
rk887 n36__i12__net2 n37__i12__net2 18.9968
rk888 n37__i12__net2 n36__i12__net2 4.4072
rk889 n7__i12__net1 n8__i12__net1 6.7179
rk890 n8__i12__net1 n9__i12__net1 15.4738
rk891 n8__i12__net1 n10__i12__net1 301.9e-3
rk892 n10__i12__net1 n4__i12__net1 45.1782
rk893 i12__net1 n10__i12__net1 45
rk895 n11__vddio n12__vddio 491.5e-3
rk896 n12__vddio n14__vddio 8.648e-3
rk897 n14__vddio n8__vddio 790e-3
rk898 n11__vddio n16__vddio 489.8e-3
rk899 n16__vddio n17__vddio 1.4774
rk900 n17__vddio n18__vddio 1.5153
rk901 n18__vddio n19__vddio 1.0928
rk902 n19__vddio n15__vddio 3.6646
rk903 n12__vddio n20__vddio 22.22e-3
rk904 n20__vddio n22__vddio 2.3235
rk905 n22__vddio n23__vddio 1.0607
rk906 n23__vddio n21__vddio 4.6153
rk907 n14__vddio n24__vddio 700.8e-3
rk908 n20__vddio n25__vddio 11.6593
rk909 n13__vddio n14__vddio 2.0833
rk910 n15__vddio n16__vddio 3.2632
rk911 n15__vddio n17__vddio 3.1
rk912 n15__vddio n18__vddio 3.1
rk913 n21__vddio n22__vddio 7.75
rk914 n21__vddio n23__vddio 3.1
rk916 n259__vss n260__vss 14.08e-3
rk917 n260__vss n261__vss 1.4701
rk918 n261__vss n262__vss 562e-3
rk919 n262__vss n263__vss 494e-3
rk920 n263__vss n264__vss 7.676e-3
rk921 n264__vss n256__vss 598.4e-3
rk923 n263__vss n266__vss 17.85e-3
rk924 n266__vss n267__vss 17.7476
rk925 n264__vss n268__vss 855.1e-3
rk926 n266__vss n270__vss 1.6452
rk927 n270__vss n269__vss 19.6592
rk928 n258__vss n259__vss 3.9474
rk929 n258__vss n261__vss 3.75
rk930 n7__vss n264__vss 1.7222
rk931 n269__vss n270__vss 3.75
rk932 n10__i12__net3 n11__i12__net3 4.7406
rk933 n11__i12__net3 n12__i12__net3 1.5153
rk934 n12__i12__net3 n13__i12__net3 1.4995
rk935 n13__i12__net3 n14__i12__net3 174.2e-3
rk937 n10__i12__net3 n11__i12__net3 3.1
rk938 n10__i12__net3 n12__i12__net3 3.1
rk939 n10__i12__net3 n13__i12__net3 3.2632
rk941 n17__i12__net3 n19__i12__net3 369.9e-3
rk942 n19__i12__net3 n18__i12__net3 5.2385
rk943 n18__i12__net3 n19__i12__net3 3.9474
rk944 n26__vddio n27__vddio 4.7406
rk945 n27__vddio n28__vddio 1.5153
rk946 n28__vddio n29__vddio 1.091
rk947 n29__vddio n26__vddio 3.6628
rk948 n26__vddio n27__vddio 3.1
rk949 n26__vddio n28__vddio 3.1
rk951 n273__vss n274__vss 14.08e-3
rk952 n274__vss n272__vss 5.2201
rk953 n272__vss n273__vss 3.9474
rk954 n26__i12__net3 n27__i12__net3 4.7406
rk955 n27__i12__net3 n28__i12__net3 1.5153
rk956 n28__i12__net3 n29__i12__net3 1.4995
rk957 n29__i12__net3 n30__i12__net3 180.5e-3
rk959 n26__i12__net3 n27__i12__net3 3.1
rk960 n26__i12__net3 n28__i12__net3 3.1
rk961 n26__i12__net3 n29__i12__net3 3.2632
rk963 n33__i12__net3 n35__i12__net3 363.6e-3
rk964 n35__i12__net3 n34__i12__net3 5.2385
rk965 n34__i12__net3 n35__i12__net3 3.9474
rk966 n30__vddio n31__vddio 4.7406
rk967 n31__vddio n32__vddio 1.5153
rk968 n32__vddio n33__vddio 1.0865
rk969 n33__vddio n30__vddio 3.6709
rk970 n30__vddio n31__vddio 3.1
rk971 n30__vddio n32__vddio 3.1
rk973 n277__vss n278__vss 8.446e-3
rk974 n278__vss n276__vss 5.2264
rk975 n276__vss n277__vss 3.9474
rk976 n42__i12__net3 n43__i12__net3 4.7406
rk977 n43__i12__net3 n44__i12__net3 1.5153
rk978 n44__i12__net3 n45__i12__net3 1.4995
rk979 n45__i12__net3 n46__i12__net3 174.2e-3
rk981 n42__i12__net3 n43__i12__net3 3.1
rk982 n42__i12__net3 n44__i12__net3 3.1
rk983 n42__i12__net3 n45__i12__net3 3.2632
rk985 n49__i12__net3 n51__i12__net3 369.9e-3
rk986 n51__i12__net3 n50__i12__net3 5.2385
rk987 n50__i12__net3 n51__i12__net3 3.9474
rk988 n34__vddio n35__vddio 4.7406
rk989 n35__vddio n36__vddio 1.5153
rk990 n36__vddio n37__vddio 1.0928
rk991 n37__vddio n34__vddio 3.6646
rk992 n34__vddio n35__vddio 3.1
rk993 n34__vddio n36__vddio 3.1
rk995 n281__vss n282__vss 14.08e-3
rk996 n282__vss n280__vss 5.2201
rk997 n280__vss n281__vss 3.9474
rk998 n58__i12__net3 n59__i12__net3 4.7406
rk999 n59__i12__net3 n60__i12__net3 1.5153
rk1000 n60__i12__net3 n61__i12__net3 1.4995
rk1001 n61__i12__net3 n62__i12__net3 180.5e-3
rk1003 n58__i12__net3 n59__i12__net3 3.1
rk1004 n58__i12__net3 n60__i12__net3 3.1
rk1005 n58__i12__net3 n61__i12__net3 3.2632
rk1007 n65__i12__net3 n67__i12__net3 363.6e-3
rk1008 n67__i12__net3 n66__i12__net3 5.2385
rk1009 n66__i12__net3 n67__i12__net3 3.9474
rk1010 n38__vddio n39__vddio 4.7406
rk1011 n39__vddio n40__vddio 1.5153
rk1012 n40__vddio n41__vddio 1.0879
rk1013 n41__vddio n38__vddio 3.666
rk1014 n38__vddio n39__vddio 3.1
rk1015 n38__vddio n40__vddio 3.1
rk1017 n285__vss n286__vss 11.26e-3
rk1018 n286__vss n284__vss 5.2233
rk1019 n284__vss n285__vss 3.9474
rk1020 n74__i12__net3 n75__i12__net3 4.7406
rk1021 n75__i12__net3 n76__i12__net3 1.5153
rk1022 n76__i12__net3 n77__i12__net3 1.4995
rk1023 n77__i12__net3 n78__i12__net3 177.3e-3
rk1025 n74__i12__net3 n75__i12__net3 3.1
rk1026 n74__i12__net3 n76__i12__net3 3.1
rk1027 n74__i12__net3 n77__i12__net3 3.2632
rk1029 n81__i12__net3 n83__i12__net3 366.7e-3
rk1030 n83__i12__net3 n82__i12__net3 5.2385
rk1031 n82__i12__net3 n83__i12__net3 3.9474
rk1032 n42__vddio n43__vddio 4.7406
rk1033 n43__vddio n44__vddio 1.5153
rk1034 n44__vddio n45__vddio 1.0928
rk1035 n45__vddio n42__vddio 3.6646
rk1036 n42__vddio n43__vddio 3.1
rk1037 n42__vddio n44__vddio 3.1
rk1039 n289__vss n290__vss 14.08e-3
rk1040 n290__vss n288__vss 5.2201
rk1041 n288__vss n289__vss 3.9474
rk1042 n43__i12__net2 n44__i12__net2 8.8107
rk1043 n44__i12__net2 n45__i12__net2 1.5153
rk1044 n45__i12__net2 n41__i12__net2 522.8e-3
rk1045 n41__i12__net2 n46__i12__net2 344e-3
rk1046 n46__i12__net2 n48__i12__net2 421.1e-3
rk1047 n48__i12__net2 n42__i12__net2 245e-3
rk1048 n42__i12__net2 n47__i12__net2 4.4054
rk1049 n46__i12__net2 n49__i12__net2 301.9e-3
rk1050 n49__i12__net2 n50__i12__net2 178.2e-3
rk1051 n50__i12__net2 n51__i12__net2 178.2e-3
rk1052 n51__i12__net2 n52__i12__net2 178.2e-3
rk1053 n52__i12__net2 n53__i12__net2 178.2e-3
rk1054 n53__i12__net2 n54__i12__net2 178.2e-3
rk1055 n54__i12__net2 n55__i12__net2 178.2e-3
rk1056 n55__i12__net2 n56__i12__net2 178.2e-3
rk1057 n56__i12__net2 n57__i12__net2 178.2e-3
rk1058 n57__i12__net2 n58__i12__net2 178.2e-3
rk1059 n58__i12__net2 n38__i12__net2 45.1782
rk1060 n43__i12__net2 n44__i12__net2 3.1
rk1061 n43__i12__net2 n45__i12__net2 3.1
rk1062 n47__i12__net2 n48__i12__net2 18.75
rk1063 i12__net2 n49__i12__net2 45
rk1064 n4__i12__net2 n50__i12__net2 45
rk1065 n7__i12__net2 n51__i12__net2 45
rk1066 n10__i12__net2 n52__i12__net2 45
rk1067 n13__i12__net2 n53__i12__net2 45
rk1068 n16__i12__net2 n54__i12__net2 45
rk1069 n19__i12__net2 n55__i12__net2 45
rk1070 n22__i12__net2 n56__i12__net2 45
rk1071 n25__i12__net2 n57__i12__net2 45
rk1072 n28__i12__net2 n58__i12__net2 45
rk1073 n1__r_out n2__r_out 4.884
rk1074 n2__r_out n3__r_out 1.5153
rk1075 n3__r_out n4__r_out 602.2e-3
rk1076 n4__r_out n1__r_out 4.1652
rk1077 n1__r_out n2__r_out 3.1
rk1078 n1__r_out n3__r_out 3.1
rk1080 n6__r_out n8__r_out 397e-3
rk1081 n8__r_out n7__r_out 5.4217
rk1082 n7__r_out n8__r_out 3.9474
rk1083 n50__vddio n51__vddio 4.884
rk1084 n51__vddio n52__vddio 1.0076
rk1085 n52__vddio n53__vddio 502.5e-3
rk1086 n53__vddio n50__vddio 4.769
rk1087 n50__vddio n51__vddio 3.1
rk1088 n50__vddio n53__vddio 3.1
rk1089 n295__vss n296__vss 4.4467
rk1090 n296__vss n295__vss 4.9171
rk1091 n9__r_out n10__r_out 4.884
rk1092 n10__r_out n11__r_out 1.5153
rk1093 n11__r_out n12__r_out 603.5e-3
rk1094 n12__r_out n9__r_out 4.1603
rk1095 n9__r_out n10__r_out 3.1
rk1096 n9__r_out n11__r_out 3.1
rk1098 n14__r_out n16__r_out 392e-3
rk1099 n16__r_out n15__r_out 5.4217
rk1100 n15__r_out n16__r_out 3.9474
rk1101 n54__vddio n55__vddio 4.884
rk1102 n55__vddio n56__vddio 1.0108
rk1103 n56__vddio n57__vddio 499.3e-3
rk1104 n57__vddio n54__vddio 4.769
rk1105 n54__vddio n55__vddio 3.1
rk1106 n54__vddio n57__vddio 3.1
rk1107 n297__vss n298__vss 4.4499
rk1108 n298__vss n297__vss 4.9139
rk1109 n17__r_out n18__r_out 4.884
rk1110 n18__r_out n19__r_out 1.5153
rk1111 n19__r_out n20__r_out 602.2e-3
rk1112 n20__r_out n17__r_out 4.1652
rk1113 n17__r_out n18__r_out 3.1
rk1114 n17__r_out n19__r_out 3.1
rk1116 n22__r_out n24__r_out 397e-3
rk1117 n24__r_out n23__r_out 5.4217
rk1118 n23__r_out n24__r_out 3.9474
rk1119 n58__vddio n59__vddio 4.884
rk1120 n59__vddio n60__vddio 1.0094
rk1121 n60__vddio n61__vddio 504.3e-3
rk1122 n61__vddio n58__vddio 4.769
rk1123 n58__vddio n59__vddio 3.1
rk1124 n58__vddio n61__vddio 3.1
rk1125 n299__vss n300__vss 4.4485
rk1126 n300__vss n299__vss 4.9189
rk1127 n25__r_out n26__r_out 4.884
rk1128 n26__r_out n27__r_out 1.5153
rk1129 n27__r_out n28__r_out 600.4e-3
rk1130 n28__r_out n25__r_out 4.1634
rk1131 n25__r_out n26__r_out 3.1
rk1132 n25__r_out n27__r_out 3.1
rk1134 n30__r_out n32__r_out 395.2e-3
rk1135 n32__r_out n31__r_out 5.4217
rk1136 n31__r_out n32__r_out 3.9474
rk1137 n62__vddio n63__vddio 4.884
rk1138 n63__vddio n64__vddio 1.0076
rk1139 n64__vddio n65__vddio 502.5e-3
rk1140 n65__vddio n62__vddio 4.769
rk1141 n62__vddio n63__vddio 3.1
rk1142 n62__vddio n65__vddio 3.1
rk1143 n301__vss n302__vss 4.4467
rk1144 n302__vss n301__vss 4.9171
rk1145 n33__r_out n34__r_out 4.884
rk1146 n34__r_out n35__r_out 1.5153
rk1147 n35__r_out n36__r_out 598.5e-3
rk1148 n36__r_out n33__r_out 4.1616
rk1149 n33__r_out n34__r_out 3.1
rk1150 n33__r_out n35__r_out 3.1
rk1152 n38__r_out n40__r_out 393.3e-3
rk1153 n40__r_out n39__r_out 5.4217
rk1154 n39__r_out n40__r_out 3.9474
rk1155 n66__vddio n67__vddio 4.884
rk1156 n67__vddio n68__vddio 1.0058
rk1157 n68__vddio n69__vddio 500.7e-3
rk1158 n69__vddio n66__vddio 4.769
rk1159 n66__vddio n67__vddio 3.1
rk1160 n66__vddio n69__vddio 3.1
rk1161 n303__vss n304__vss 4.4449
rk1162 n304__vss n303__vss 4.9153
rk1163 n41__r_out n42__r_out 4.884
rk1164 n42__r_out n43__r_out 1.5153
rk1165 n43__r_out n44__r_out 603.5e-3
rk1166 n44__r_out n41__r_out 4.1603
rk1167 n41__r_out n42__r_out 3.1
rk1168 n41__r_out n43__r_out 3.1
rk1170 n46__r_out n48__r_out 392e-3
rk1171 n48__r_out n47__r_out 5.4217
rk1172 n47__r_out n48__r_out 3.9474
rk1173 n70__vddio n71__vddio 4.884
rk1174 n71__vddio n72__vddio 1.0108
rk1175 n72__vddio n73__vddio 499.3e-3
rk1176 n73__vddio n70__vddio 4.769
rk1177 n70__vddio n71__vddio 3.1
rk1178 n70__vddio n73__vddio 3.1
rk1179 n305__vss n306__vss 4.4499
rk1180 n306__vss n305__vss 4.9139
rk1181 n49__r_out n50__r_out 4.884
rk1182 n50__r_out n51__r_out 1.5153
rk1183 n51__r_out n52__r_out 600.4e-3
rk1184 n52__r_out n49__r_out 4.1634
rk1185 n49__r_out n50__r_out 3.1
rk1186 n49__r_out n51__r_out 3.1
rk1188 n54__r_out n56__r_out 395.2e-3
rk1189 n56__r_out n55__r_out 5.4217
rk1190 n55__r_out n56__r_out 3.9474
rk1191 n74__vddio n75__vddio 4.884
rk1192 n75__vddio n76__vddio 1.0076
rk1193 n76__vddio n77__vddio 502.5e-3
rk1194 n77__vddio n74__vddio 4.769
rk1195 n74__vddio n75__vddio 3.1
rk1196 n74__vddio n77__vddio 3.1
rk1197 n307__vss n308__vss 4.4467
rk1198 n308__vss n307__vss 4.9171
rk1199 n57__r_out n58__r_out 4.884
rk1200 n58__r_out n59__r_out 1.5153
rk1201 n59__r_out n60__r_out 598.5e-3
rk1202 n60__r_out n57__r_out 4.1616
rk1203 n57__r_out n58__r_out 3.1
rk1204 n57__r_out n59__r_out 3.1
rk1206 n62__r_out n64__r_out 393.3e-3
rk1207 n64__r_out n63__r_out 5.4217
rk1208 n63__r_out n64__r_out 3.9474
rk1209 n78__vddio n79__vddio 4.884
rk1210 n79__vddio n80__vddio 1.0058
rk1211 n80__vddio n81__vddio 500.7e-3
rk1212 n81__vddio n78__vddio 4.769
rk1213 n78__vddio n79__vddio 3.1
rk1214 n78__vddio n81__vddio 3.1
rk1215 n309__vss n310__vss 4.4449
rk1216 n310__vss n309__vss 4.9153
rk1217 n65__r_out n66__r_out 4.884
rk1218 n66__r_out n67__r_out 1.5153
rk1219 n67__r_out n68__r_out 603.5e-3
rk1220 n68__r_out n65__r_out 4.1603
rk1221 n65__r_out n66__r_out 3.1
rk1222 n65__r_out n67__r_out 3.1
rk1224 n70__r_out n72__r_out 392e-3
rk1225 n72__r_out n71__r_out 5.4217
rk1226 n71__r_out n72__r_out 3.9474
rk1227 n82__vddio n83__vddio 4.884
rk1228 n83__vddio n84__vddio 1.0108
rk1229 n84__vddio n85__vddio 499.3e-3
rk1230 n85__vddio n82__vddio 4.769
rk1231 n82__vddio n83__vddio 3.1
rk1232 n82__vddio n85__vddio 3.1
rk1233 n311__vss n312__vss 4.4499
rk1234 n312__vss n311__vss 4.9139
rk1235 n73__r_out n74__r_out 4.884
rk1236 n74__r_out n75__r_out 1.5153
rk1237 n75__r_out n76__r_out 600.4e-3
rk1238 n76__r_out n73__r_out 4.1634
rk1239 n73__r_out n74__r_out 3.1
rk1240 n73__r_out n75__r_out 3.1
rk1242 n78__r_out n80__r_out 395.2e-3
rk1243 n80__r_out n79__r_out 5.4217
rk1244 n79__r_out n80__r_out 3.9474
rk1245 n86__vddio n87__vddio 4.884
rk1246 n87__vddio n88__vddio 1.0076
rk1247 n88__vddio n89__vddio 502.5e-3
rk1248 n89__vddio n86__vddio 4.769
rk1249 n86__vddio n87__vddio 3.1
rk1250 n86__vddio n89__vddio 3.1
rk1251 n313__vss n314__vss 4.4467
rk1252 n314__vss n313__vss 4.9171
rk1253 n81__r_out n82__r_out 4.884
rk1254 n82__r_out n83__r_out 1.5153
rk1255 n83__r_out n84__r_out 602.4e-3
rk1256 n84__r_out n81__r_out 4.1655
rk1257 n81__r_out n82__r_out 3.1
rk1258 n81__r_out n83__r_out 3.1
rk1260 n86__r_out n88__r_out 397.2e-3
rk1261 n88__r_out n87__r_out 5.4217
rk1262 n87__r_out n88__r_out 3.9474
rk1263 n90__vddio n91__vddio 4.884
rk1264 n91__vddio n92__vddio 1.0097
rk1265 n92__vddio n93__vddio 504.6e-3
rk1266 n93__vddio n90__vddio 4.769
rk1267 n90__vddio n91__vddio 3.1
rk1268 n90__vddio n93__vddio 3.1
rk1269 n315__vss n316__vss 4.4488
rk1270 n316__vss n315__vss 4.9192
rk1271 n89__r_out n90__r_out 4.884
rk1272 n90__r_out n91__r_out 1.5153
rk1273 n91__r_out n92__r_out 605.3e-3
rk1274 n92__r_out n89__r_out 4.1621
rk1275 n89__r_out n90__r_out 3.1
rk1276 n89__r_out n91__r_out 3.1
rk1278 n94__r_out n96__r_out 393.8e-3
rk1279 n96__r_out n95__r_out 5.4217
rk1280 n95__r_out n96__r_out 3.9474
rk1281 n94__vddio n95__vddio 4.884
rk1282 n95__vddio n96__vddio 1.0126
rk1283 n96__vddio n97__vddio 501.2e-3
rk1284 n97__vddio n94__vddio 4.769
rk1285 n94__vddio n95__vddio 3.1
rk1286 n94__vddio n97__vddio 3.1
rk1287 n317__vss n318__vss 4.4517
rk1288 n318__vss n317__vss 4.9158
rk1289 n97__r_out n98__r_out 4.884
rk1290 n98__r_out n99__r_out 1.5153
rk1291 n99__r_out n100__r_out 598.5e-3
rk1292 n100__r_out n97__r_out 4.1616
rk1293 n97__r_out n98__r_out 3.1
rk1294 n97__r_out n99__r_out 3.1
rk1296 n102__r_out n104__r_out 393.3e-3
rk1297 n104__r_out n103__r_out 5.4217
rk1298 n103__r_out n104__r_out 3.9474
rk1299 n98__vddio n99__vddio 4.884
rk1300 n99__vddio n100__vddio 1.0058
rk1301 n100__vddio n101__vddio 500.7e-3
rk1302 n101__vddio n98__vddio 4.769
rk1303 n98__vddio n99__vddio 3.1
rk1304 n98__vddio n101__vddio 3.1
rk1305 n319__vss n320__vss 4.4449
rk1306 n320__vss n319__vss 4.9153
rk1307 n105__r_out n106__r_out 4.884
rk1308 n106__r_out n107__r_out 1.5153
rk1309 n107__r_out n108__r_out 602.4e-3
rk1310 n108__r_out n105__r_out 4.1655
rk1311 n105__r_out n106__r_out 3.1
rk1312 n105__r_out n107__r_out 3.1
rk1314 n110__r_out n112__r_out 397.2e-3
rk1315 n112__r_out n111__r_out 5.4217
rk1316 n111__r_out n112__r_out 3.9474
rk1317 n102__vddio n103__vddio 4.884
rk1318 n103__vddio n104__vddio 1.0097
rk1319 n104__vddio n105__vddio 504.6e-3
rk1320 n105__vddio n102__vddio 4.769
rk1321 n102__vddio n103__vddio 3.1
rk1322 n102__vddio n105__vddio 3.1
rk1323 n321__vss n322__vss 4.4488
rk1324 n322__vss n321__vss 4.9192
rk1325 n113__r_out n114__r_out 4.884
rk1326 n114__r_out n115__r_out 1.5153
rk1327 n115__r_out n116__r_out 605.3e-3
rk1328 n116__r_out n113__r_out 4.1621
rk1329 n113__r_out n114__r_out 3.1
rk1330 n113__r_out n115__r_out 3.1
rk1332 n118__r_out n120__r_out 393.8e-3
rk1333 n120__r_out n119__r_out 5.4217
rk1334 n119__r_out n120__r_out 3.9474
rk1335 n106__vddio n107__vddio 4.884
rk1336 n107__vddio n108__vddio 1.0126
rk1337 n108__vddio n109__vddio 501.2e-3
rk1338 n109__vddio n106__vddio 4.769
rk1339 n106__vddio n107__vddio 3.1
rk1340 n106__vddio n109__vddio 3.1
rk1341 n323__vss n324__vss 4.4517
rk1342 n324__vss n323__vss 4.9158
rk1343 n121__r_out n122__r_out 4.884
rk1344 n122__r_out n123__r_out 1.5153
rk1345 n123__r_out n124__r_out 598.5e-3
rk1346 n124__r_out n121__r_out 4.1616
rk1347 n121__r_out n122__r_out 3.1
rk1348 n121__r_out n123__r_out 3.1
rk1350 n126__r_out n128__r_out 393.3e-3
rk1351 n128__r_out n127__r_out 5.4217
rk1352 n127__r_out n128__r_out 3.9474
rk1353 n110__vddio n111__vddio 4.884
rk1354 n111__vddio n112__vddio 1.0058
rk1355 n112__vddio n113__vddio 500.7e-3
rk1356 n113__vddio n110__vddio 4.769
rk1357 n110__vddio n111__vddio 3.1
rk1358 n110__vddio n113__vddio 3.1
rk1359 n325__vss n326__vss 4.4449
rk1360 n326__vss n325__vss 4.9153
rk1361 n129__r_out n130__r_out 4.884
rk1362 n130__r_out n131__r_out 1.5153
rk1363 n131__r_out n132__r_out 600.4e-3
rk1364 n132__r_out n129__r_out 4.1634
rk1365 n129__r_out n130__r_out 3.1
rk1366 n129__r_out n131__r_out 3.1
rk1368 n134__r_out n136__r_out 395.2e-3
rk1369 n136__r_out n135__r_out 5.4217
rk1370 n135__r_out n136__r_out 3.9474
rk1371 n114__vddio n115__vddio 4.884
rk1372 n115__vddio n116__vddio 1.0076
rk1373 n116__vddio n117__vddio 502.5e-3
rk1374 n117__vddio n114__vddio 4.769
rk1375 n114__vddio n115__vddio 3.1
rk1376 n114__vddio n117__vddio 3.1
rk1377 n327__vss n328__vss 4.4467
rk1378 n328__vss n327__vss 4.9171
rk1379 n137__r_out n138__r_out 4.884
rk1380 n138__r_out n139__r_out 1.5153
rk1381 n139__r_out n140__r_out 603.5e-3
rk1382 n140__r_out n137__r_out 4.1603
rk1383 n137__r_out n138__r_out 3.1
rk1384 n137__r_out n139__r_out 3.1
rk1386 n142__r_out n144__r_out 392e-3
rk1387 n144__r_out n143__r_out 5.4217
rk1388 n143__r_out n144__r_out 3.9474
rk1389 n118__vddio n119__vddio 4.884
rk1390 n119__vddio n120__vddio 1.0108
rk1391 n120__vddio n121__vddio 499.3e-3
rk1392 n121__vddio n118__vddio 4.769
rk1393 n118__vddio n119__vddio 3.1
rk1394 n118__vddio n121__vddio 3.1
rk1395 n329__vss n330__vss 4.4499
rk1396 n330__vss n329__vss 4.9139
rk1397 n145__r_out n146__r_out 4.884
rk1398 n146__r_out n147__r_out 1.5153
rk1399 n147__r_out n148__r_out 602.2e-3
rk1400 n148__r_out n145__r_out 4.1652
rk1401 n145__r_out n146__r_out 3.1
rk1402 n145__r_out n147__r_out 3.1
rk1404 n150__r_out n152__r_out 397e-3
rk1405 n152__r_out n151__r_out 5.4217
rk1406 n151__r_out n152__r_out 3.9474
rk1407 n122__vddio n123__vddio 4.884
rk1408 n123__vddio n124__vddio 1.0094
rk1409 n124__vddio n125__vddio 504.3e-3
rk1410 n125__vddio n122__vddio 4.769
rk1411 n122__vddio n123__vddio 3.1
rk1412 n122__vddio n125__vddio 3.1
rk1413 n331__vss n332__vss 4.4485
rk1414 n332__vss n331__vss 4.9189
rk1415 n153__r_out n154__r_out 4.884
rk1416 n154__r_out n155__r_out 1.5153
rk1417 n155__r_out n156__r_out 600.4e-3
rk1418 n156__r_out n153__r_out 4.1634
rk1419 n153__r_out n154__r_out 3.1
rk1420 n153__r_out n155__r_out 3.1
rk1422 n158__r_out n160__r_out 395.2e-3
rk1423 n160__r_out n159__r_out 5.4217
rk1424 n159__r_out n160__r_out 3.9474
rk1425 n126__vddio n127__vddio 4.884
rk1426 n127__vddio n128__vddio 1.0076
rk1427 n128__vddio n129__vddio 502.5e-3
rk1428 n129__vddio n126__vddio 4.769
rk1429 n126__vddio n127__vddio 3.1
rk1430 n126__vddio n129__vddio 3.1
rk1431 n333__vss n334__vss 4.4467
rk1432 n334__vss n333__vss 4.9171
rk1433 n161__r_out n162__r_out 4.884
rk1434 n162__r_out n163__r_out 1.5153
rk1435 n163__r_out n164__r_out 603.5e-3
rk1436 n164__r_out n161__r_out 4.1603
rk1437 n161__r_out n162__r_out 3.1
rk1438 n161__r_out n163__r_out 3.1
rk1440 n166__r_out n168__r_out 392e-3
rk1441 n168__r_out n167__r_out 5.4217
rk1442 n167__r_out n168__r_out 3.9474
rk1443 n130__vddio n131__vddio 4.884
rk1444 n131__vddio n132__vddio 1.0108
rk1445 n132__vddio n133__vddio 499.3e-3
rk1446 n133__vddio n130__vddio 4.769
rk1447 n130__vddio n131__vddio 3.1
rk1448 n130__vddio n133__vddio 3.1
rk1449 n335__vss n336__vss 4.4499
rk1450 n336__vss n335__vss 4.9139
rk1451 n169__r_out n170__r_out 4.884
rk1452 n170__r_out n171__r_out 1.5153
rk1453 n171__r_out n172__r_out 602.2e-3
rk1454 n172__r_out n169__r_out 4.1652
rk1455 n169__r_out n170__r_out 3.1
rk1456 n169__r_out n171__r_out 3.1
rk1458 n174__r_out n176__r_out 397e-3
rk1459 n176__r_out n175__r_out 5.4217
rk1460 n175__r_out n176__r_out 3.9474
rk1461 n135__vddio n136__vddio 504.3e-3
rk1462 n136__vddio n137__vddio 1.0094
rk1463 n137__vddio n138__vddio 1.4396
rk1464 n138__vddio n13__vddio 25.8778
rk1465 n135__vddio n134__vddio 4.769
rk1466 n134__vddio n135__vddio 3.1
rk1467 n134__vddio n137__vddio 3.1
rk1468 n134__vddio n138__vddio 3.4444
rk1469 n337__vss n338__vss 4.4485
rk1470 n338__vss n339__vss 971.5e-3
rk1471 n339__vss n7__vss 7.8279
rk1472 n337__vss n339__vss 3.9474
rk1474 n178__r_out n180__r_out 395.2e-3
rk1475 n180__r_out n179__r_out 5.4217
rk1476 n179__r_out n180__r_out 3.9474
rk1477 n181__r_out n182__r_out 4.884
rk1478 n182__r_out n183__r_out 1.5153
rk1479 n183__r_out n184__r_out 602.2e-3
rk1480 n184__r_out n181__r_out 4.1652
rk1481 n181__r_out n182__r_out 3.1
rk1482 n181__r_out n183__r_out 3.1
rk1483 n139__vddio n140__vddio 4.884
rk1484 n140__vddio n141__vddio 1.0076
rk1485 n141__vddio n142__vddio 502.5e-3
rk1486 n142__vddio n139__vddio 4.769
rk1487 n139__vddio n140__vddio 3.1
rk1488 n139__vddio n142__vddio 3.1
rk1489 n340__vss n341__vss 4.4467
rk1490 n341__vss n340__vss 4.9171
rk1491 n185__r_out n186__r_out 4.884
rk1492 n186__r_out n187__r_out 1.5153
rk1493 n187__r_out n188__r_out 603.5e-3
rk1494 n188__r_out n185__r_out 4.1603
rk1495 n185__r_out n186__r_out 3.1
rk1496 n185__r_out n187__r_out 3.1
rk1498 n190__r_out n192__r_out 392e-3
rk1499 n192__r_out n191__r_out 5.4217
rk1500 n191__r_out n192__r_out 3.9474
rk1501 n143__vddio n144__vddio 4.884
rk1502 n144__vddio n145__vddio 1.0108
rk1503 n145__vddio n146__vddio 499.3e-3
rk1504 n146__vddio n143__vddio 4.769
rk1505 n143__vddio n144__vddio 3.1
rk1506 n143__vddio n146__vddio 3.1
rk1507 n342__vss n343__vss 4.4499
rk1508 n343__vss n342__vss 4.9139
rk1509 n193__r_out n194__r_out 4.884
rk1510 n194__r_out n195__r_out 1.5153
rk1511 n195__r_out n196__r_out 602.2e-3
rk1512 n196__r_out n193__r_out 4.1652
rk1513 n193__r_out n194__r_out 3.1
rk1514 n193__r_out n195__r_out 3.1
rk1516 n198__r_out n200__r_out 397e-3
rk1517 n200__r_out n199__r_out 5.4217
rk1518 n199__r_out n200__r_out 3.9474
rk1519 n147__vddio n148__vddio 4.884
rk1520 n148__vddio n149__vddio 1.0094
rk1521 n149__vddio n150__vddio 504.3e-3
rk1522 n150__vddio n147__vddio 4.769
rk1523 n147__vddio n148__vddio 3.1
rk1524 n147__vddio n150__vddio 3.1
rk1525 n344__vss n345__vss 4.4485
rk1526 n345__vss n344__vss 4.9189
rk1527 n201__r_out n202__r_out 4.884
rk1528 n202__r_out n203__r_out 1.5153
rk1529 n203__r_out n204__r_out 600.4e-3
rk1530 n204__r_out n201__r_out 4.1634
rk1531 n201__r_out n202__r_out 3.1
rk1532 n201__r_out n203__r_out 3.1
rk1534 n206__r_out n208__r_out 395.2e-3
rk1535 n208__r_out n207__r_out 5.4217
rk1536 n207__r_out n208__r_out 3.9474
rk1537 n151__vddio n152__vddio 4.884
rk1538 n152__vddio n153__vddio 1.0076
rk1539 n153__vddio n154__vddio 502.5e-3
rk1540 n154__vddio n151__vddio 4.769
rk1541 n151__vddio n152__vddio 3.1
rk1542 n151__vddio n154__vddio 3.1
rk1543 n346__vss n347__vss 4.4467
rk1544 n347__vss n346__vss 4.9171
rk1545 n209__r_out n210__r_out 4.884
rk1546 n210__r_out n211__r_out 1.5153
rk1547 n211__r_out n212__r_out 603.5e-3
rk1548 n212__r_out n209__r_out 4.1603
rk1549 n209__r_out n210__r_out 3.1
rk1550 n209__r_out n211__r_out 3.1
rk1552 n214__r_out n216__r_out 392e-3
rk1553 n216__r_out n215__r_out 5.4217
rk1554 n215__r_out n216__r_out 3.9474
rk1555 n155__vddio n156__vddio 4.884
rk1556 n156__vddio n157__vddio 1.0108
rk1557 n157__vddio n158__vddio 499.3e-3
rk1558 n158__vddio n155__vddio 4.769
rk1559 n155__vddio n156__vddio 3.1
rk1560 n155__vddio n158__vddio 3.1
rk1561 n348__vss n349__vss 4.4499
rk1562 n349__vss n348__vss 4.9139
rk1563 n217__r_out n218__r_out 4.884
rk1564 n218__r_out n219__r_out 1.5153
rk1565 n219__r_out n220__r_out 602.9e-3
rk1566 n220__r_out n217__r_out 4.166
rk1567 n217__r_out n218__r_out 3.1
rk1568 n217__r_out n219__r_out 3.1
rk1570 n222__r_out n224__r_out 397.7e-3
rk1571 n224__r_out n223__r_out 5.4217
rk1572 n223__r_out n224__r_out 3.9474
rk1573 n159__vddio n160__vddio 4.884
rk1574 n160__vddio n161__vddio 1.0102
rk1575 n161__vddio n162__vddio 505e-3
rk1576 n162__vddio n159__vddio 4.769
rk1577 n159__vddio n160__vddio 3.1
rk1578 n159__vddio n162__vddio 3.1
rk1579 n350__vss n351__vss 4.4493
rk1580 n351__vss n350__vss 4.9196
rk1581 n225__r_out n226__r_out 4.884
rk1582 n226__r_out n227__r_out 1.5153
rk1583 n227__r_out n228__r_out 605.6e-3
rk1584 n228__r_out n225__r_out 4.1624
rk1585 n225__r_out n226__r_out 3.1
rk1586 n225__r_out n227__r_out 3.1
rk1588 n230__r_out n232__r_out 394.1e-3
rk1589 n232__r_out n231__r_out 5.4217
rk1590 n231__r_out n232__r_out 3.9474
rk1591 n163__vddio n164__vddio 4.884
rk1592 n164__vddio n165__vddio 1.0128
rk1593 n165__vddio n166__vddio 501.4e-3
rk1594 n166__vddio n163__vddio 4.769
rk1595 n163__vddio n164__vddio 3.1
rk1596 n163__vddio n166__vddio 3.1
rk1597 n352__vss n353__vss 4.4519
rk1598 n353__vss n352__vss 4.916
rk1599 n233__r_out n234__r_out 4.884
rk1600 n234__r_out n235__r_out 1.5153
rk1601 n235__r_out n236__r_out 602.2e-3
rk1602 n236__r_out n233__r_out 4.1652
rk1603 n233__r_out n234__r_out 3.1
rk1604 n233__r_out n235__r_out 3.1
rk1606 n238__r_out n240__r_out 397e-3
rk1607 n240__r_out n239__r_out 5.4217
rk1608 n239__r_out n240__r_out 3.9474
rk1609 n167__vddio n168__vddio 4.884
rk1610 n168__vddio n169__vddio 1.0094
rk1611 n169__vddio n170__vddio 504.3e-3
rk1612 n170__vddio n167__vddio 4.769
rk1613 n167__vddio n168__vddio 3.1
rk1614 n167__vddio n170__vddio 3.1
rk1615 n354__vss n355__vss 4.4485
rk1616 n355__vss n354__vss 4.9189
rk1617 n241__r_out n242__r_out 4.884
rk1618 n242__r_out n243__r_out 1.5153
rk1619 n243__r_out n244__r_out 602.9e-3
rk1620 n244__r_out n241__r_out 4.166
rk1621 n241__r_out n242__r_out 3.1
rk1622 n241__r_out n243__r_out 3.1
rk1624 n246__r_out n248__r_out 397.7e-3
rk1625 n248__r_out n247__r_out 5.4217
rk1626 n247__r_out n248__r_out 3.9474
rk1627 n171__vddio n172__vddio 4.884
rk1628 n172__vddio n173__vddio 1.0102
rk1629 n173__vddio n174__vddio 505e-3
rk1630 n174__vddio n171__vddio 4.769
rk1631 n171__vddio n172__vddio 3.1
rk1632 n171__vddio n174__vddio 3.1
rk1633 n356__vss n357__vss 4.4493
rk1634 n357__vss n356__vss 4.9196
rk1635 n249__r_out n250__r_out 4.884
rk1636 n250__r_out n251__r_out 1.5153
rk1637 n251__r_out n252__r_out 605.6e-3
rk1638 n252__r_out n249__r_out 4.1624
rk1639 n249__r_out n250__r_out 3.1
rk1640 n249__r_out n251__r_out 3.1
rk1642 n254__r_out n256__r_out 394.1e-3
rk1643 n256__r_out n255__r_out 5.4217
rk1644 n255__r_out n256__r_out 3.9474
rk1645 n175__vddio n176__vddio 4.884
rk1646 n176__vddio n177__vddio 1.0128
rk1647 n177__vddio n178__vddio 501.4e-3
rk1648 n178__vddio n175__vddio 4.769
rk1649 n175__vddio n176__vddio 3.1
rk1650 n175__vddio n178__vddio 3.1
rk1651 n358__vss n359__vss 4.4519
rk1652 n359__vss n358__vss 4.916
rk1653 n257__r_out n258__r_out 4.884
rk1654 n258__r_out n259__r_out 1.5153
rk1655 n259__r_out n260__r_out 602.2e-3
rk1656 n260__r_out n257__r_out 4.1652
rk1657 n257__r_out n258__r_out 3.1
rk1658 n257__r_out n259__r_out 3.1
rk1660 n262__r_out n264__r_out 397e-3
rk1661 n264__r_out n263__r_out 5.4217
rk1662 n263__r_out n264__r_out 3.9474
rk1663 n179__vddio n180__vddio 4.884
rk1664 n180__vddio n181__vddio 1.0094
rk1665 n181__vddio n182__vddio 504.3e-3
rk1666 n182__vddio n179__vddio 4.769
rk1667 n179__vddio n180__vddio 3.1
rk1668 n179__vddio n182__vddio 3.1
rk1669 n360__vss n361__vss 4.4485
rk1670 n361__vss n360__vss 4.9189
rk1671 n265__r_out n266__r_out 4.884
rk1672 n266__r_out n267__r_out 1.5153
rk1673 n267__r_out n268__r_out 602.9e-3
rk1674 n268__r_out n265__r_out 4.166
rk1675 n265__r_out n266__r_out 3.1
rk1676 n265__r_out n267__r_out 3.1
rk1678 n270__r_out n272__r_out 397.7e-3
rk1679 n272__r_out n271__r_out 5.4217
rk1680 n271__r_out n272__r_out 3.9474
rk1681 n183__vddio n184__vddio 4.884
rk1682 n184__vddio n185__vddio 1.0102
rk1683 n185__vddio n186__vddio 505e-3
rk1684 n186__vddio n183__vddio 4.769
rk1685 n183__vddio n184__vddio 3.1
rk1686 n183__vddio n186__vddio 3.1
rk1687 n362__vss n363__vss 4.4493
rk1688 n363__vss n362__vss 4.9196
rk1689 n273__r_out n274__r_out 4.884
rk1690 n274__r_out n275__r_out 1.5153
rk1691 n275__r_out n276__r_out 605.6e-3
rk1692 n276__r_out n273__r_out 4.1624
rk1693 n273__r_out n274__r_out 3.1
rk1694 n273__r_out n275__r_out 3.1
rk1696 n278__r_out n280__r_out 394.1e-3
rk1697 n280__r_out n279__r_out 5.4217
rk1698 n279__r_out n280__r_out 3.9474
rk1699 n187__vddio n188__vddio 4.884
rk1700 n188__vddio n189__vddio 1.0128
rk1701 n189__vddio n190__vddio 501.4e-3
rk1702 n190__vddio n187__vddio 4.769
rk1703 n187__vddio n188__vddio 3.1
rk1704 n187__vddio n190__vddio 3.1
rk1705 n364__vss n365__vss 4.4519
rk1706 n365__vss n364__vss 4.916
rk1707 n281__r_out n282__r_out 4.884
rk1708 n282__r_out n283__r_out 1.5153
rk1709 n283__r_out n284__r_out 602.2e-3
rk1710 n284__r_out n281__r_out 4.1652
rk1711 n281__r_out n282__r_out 3.1
rk1712 n281__r_out n283__r_out 3.1
rk1714 n286__r_out n288__r_out 397e-3
rk1715 n288__r_out n287__r_out 5.4217
rk1716 n287__r_out n288__r_out 3.9474
rk1717 n191__vddio n192__vddio 4.884
rk1718 n192__vddio n193__vddio 1.0094
rk1719 n193__vddio n194__vddio 504.3e-3
rk1720 n194__vddio n191__vddio 4.769
rk1721 n191__vddio n192__vddio 3.1
rk1722 n191__vddio n194__vddio 3.1
rk1723 n366__vss n367__vss 4.4485
rk1724 n367__vss n366__vss 4.9189
rk1725 n289__r_out n290__r_out 4.884
rk1726 n290__r_out n291__r_out 1.5153
rk1727 n291__r_out n292__r_out 602.9e-3
rk1728 n292__r_out n289__r_out 4.166
rk1729 n289__r_out n290__r_out 3.1
rk1730 n289__r_out n291__r_out 3.1
rk1732 n294__r_out n296__r_out 397.7e-3
rk1733 n296__r_out n295__r_out 5.4217
rk1734 n295__r_out n296__r_out 3.9474
rk1735 n195__vddio n196__vddio 4.884
rk1736 n196__vddio n197__vddio 1.0102
rk1737 n197__vddio n198__vddio 505e-3
rk1738 n198__vddio n195__vddio 4.769
rk1739 n195__vddio n196__vddio 3.1
rk1740 n195__vddio n198__vddio 3.1
rk1741 n368__vss n369__vss 4.4493
rk1742 n369__vss n368__vss 4.9196
rk1743 n297__r_out n298__r_out 4.884
rk1744 n298__r_out n299__r_out 1.5153
rk1745 n299__r_out n300__r_out 605.6e-3
rk1746 n300__r_out n297__r_out 4.1624
rk1747 n297__r_out n298__r_out 3.1
rk1748 n297__r_out n299__r_out 3.1
rk1750 n302__r_out n304__r_out 394.1e-3
rk1751 n304__r_out n303__r_out 5.4217
rk1752 n303__r_out n304__r_out 3.9474
rk1753 n199__vddio n200__vddio 4.884
rk1754 n200__vddio n201__vddio 1.0128
rk1755 n201__vddio n202__vddio 501.4e-3
rk1756 n202__vddio n199__vddio 4.769
rk1757 n199__vddio n200__vddio 3.1
rk1758 n199__vddio n202__vddio 3.1
rk1759 n370__vss n371__vss 4.4519
rk1760 n371__vss n370__vss 4.916
rk1761 n305__r_out n306__r_out 4.884
rk1762 n306__r_out n307__r_out 1.5153
rk1763 n307__r_out n308__r_out 602.2e-3
rk1764 n308__r_out n305__r_out 4.1652
rk1765 n305__r_out n306__r_out 3.1
rk1766 n305__r_out n307__r_out 3.1
rk1768 n310__r_out n312__r_out 397e-3
rk1769 n312__r_out n311__r_out 5.4217
rk1770 n311__r_out n312__r_out 3.9474
rk1771 n203__vddio n204__vddio 4.884
rk1772 n204__vddio n205__vddio 1.0094
rk1773 n205__vddio n206__vddio 504.3e-3
rk1774 n206__vddio n203__vddio 4.769
rk1775 n203__vddio n204__vddio 3.1
rk1776 n203__vddio n206__vddio 3.1
rk1777 n372__vss n373__vss 4.4485
rk1778 n373__vss n372__vss 4.9189
rk1779 n313__r_out n314__r_out 4.884
rk1780 n314__r_out n315__r_out 1.5153
rk1781 n315__r_out n316__r_out 598.5e-3
rk1782 n316__r_out n313__r_out 4.1616
rk1783 n313__r_out n314__r_out 3.1
rk1784 n313__r_out n315__r_out 3.1
rk1786 n318__r_out n320__r_out 393.3e-3
rk1787 n320__r_out n319__r_out 5.4217
rk1788 n319__r_out n320__r_out 3.9474
rk1789 n207__vddio n208__vddio 4.884
rk1790 n208__vddio n209__vddio 1.0058
rk1791 n209__vddio n210__vddio 500.7e-3
rk1792 n210__vddio n207__vddio 4.769
rk1793 n207__vddio n208__vddio 3.1
rk1794 n207__vddio n210__vddio 3.1
rk1795 n374__vss n375__vss 4.4449
rk1796 n375__vss n374__vss 4.9153
rk1797 n321__r_out n322__r_out 4.884
rk1798 n322__r_out n323__r_out 1.5153
rk1799 n323__r_out n324__r_out 603.5e-3
rk1800 n324__r_out n321__r_out 4.1603
rk1801 n321__r_out n322__r_out 3.1
rk1802 n321__r_out n323__r_out 3.1
rk1804 n326__r_out n328__r_out 392e-3
rk1805 n328__r_out n327__r_out 5.4217
rk1806 n327__r_out n328__r_out 3.9474
rk1807 n211__vddio n212__vddio 4.884
rk1808 n212__vddio n213__vddio 1.0108
rk1809 n213__vddio n214__vddio 499.3e-3
rk1810 n214__vddio n211__vddio 4.769
rk1811 n211__vddio n212__vddio 3.1
rk1812 n211__vddio n214__vddio 3.1
rk1813 n376__vss n377__vss 4.4499
rk1814 n377__vss n376__vss 4.9139
rk1815 n329__r_out n330__r_out 4.884
rk1816 n330__r_out n331__r_out 1.5153
rk1817 n331__r_out n332__r_out 600.4e-3
rk1818 n332__r_out n329__r_out 4.1634
rk1819 n329__r_out n330__r_out 3.1
rk1820 n329__r_out n331__r_out 3.1
rk1822 n334__r_out n336__r_out 395.2e-3
rk1823 n336__r_out n335__r_out 5.4217
rk1824 n335__r_out n336__r_out 3.9474
rk1825 n215__vddio n216__vddio 4.884
rk1826 n216__vddio n217__vddio 1.0076
rk1827 n217__vddio n218__vddio 502.5e-3
rk1828 n218__vddio n215__vddio 4.769
rk1829 n215__vddio n216__vddio 3.1
rk1830 n215__vddio n218__vddio 3.1
rk1831 n378__vss n379__vss 4.4467
rk1832 n379__vss n378__vss 4.9171
rk1833 n337__r_out n338__r_out 4.884
rk1834 n338__r_out n339__r_out 1.5153
rk1835 n339__r_out n340__r_out 598.5e-3
rk1836 n340__r_out n337__r_out 4.1616
rk1837 n337__r_out n338__r_out 3.1
rk1838 n337__r_out n339__r_out 3.1
rk1840 n342__r_out n344__r_out 393.3e-3
rk1841 n344__r_out n343__r_out 5.4217
rk1842 n343__r_out n344__r_out 3.9474
rk1843 n219__vddio n220__vddio 4.884
rk1844 n220__vddio n221__vddio 1.0058
rk1845 n221__vddio n222__vddio 500.7e-3
rk1846 n222__vddio n219__vddio 4.769
rk1847 n219__vddio n220__vddio 3.1
rk1848 n219__vddio n222__vddio 3.1
rk1849 n380__vss n381__vss 4.4449
rk1850 n381__vss n380__vss 4.9153
rk1851 n345__r_out n346__r_out 4.884
rk1852 n346__r_out n347__r_out 1.5153
rk1853 n347__r_out n348__r_out 603.5e-3
rk1854 n348__r_out n345__r_out 4.1603
rk1855 n345__r_out n346__r_out 3.1
rk1856 n345__r_out n347__r_out 3.1
rk1858 n350__r_out n352__r_out 392e-3
rk1859 n352__r_out n351__r_out 5.4217
rk1860 n351__r_out n352__r_out 3.9474
rk1861 n223__vddio n224__vddio 4.884
rk1862 n224__vddio n225__vddio 1.0108
rk1863 n225__vddio n226__vddio 499.3e-3
rk1864 n226__vddio n223__vddio 4.769
rk1865 n223__vddio n224__vddio 3.1
rk1866 n223__vddio n226__vddio 3.1
rk1867 n382__vss n383__vss 4.4499
rk1868 n383__vss n382__vss 4.9139
rk1869 n353__r_out n354__r_out 4.884
rk1870 n354__r_out n355__r_out 1.5153
rk1871 n355__r_out n356__r_out 600.4e-3
rk1872 n356__r_out n353__r_out 4.1634
rk1873 n353__r_out n354__r_out 3.1
rk1874 n353__r_out n355__r_out 3.1
rk1876 n358__r_out n360__r_out 395.2e-3
rk1877 n360__r_out n359__r_out 5.4217
rk1878 n359__r_out n360__r_out 3.9474
rk1879 n227__vddio n228__vddio 4.884
rk1880 n228__vddio n229__vddio 1.0076
rk1881 n229__vddio n230__vddio 502.5e-3
rk1882 n230__vddio n227__vddio 4.769
rk1883 n227__vddio n228__vddio 3.1
rk1884 n227__vddio n230__vddio 3.1
rk1885 n384__vss n385__vss 4.4467
rk1886 n385__vss n384__vss 4.9171
rk1887 n361__r_out n362__r_out 4.884
rk1888 n362__r_out n363__r_out 1.5153
rk1889 n363__r_out n364__r_out 598.5e-3
rk1890 n364__r_out n361__r_out 4.1616
rk1891 n361__r_out n362__r_out 3.1
rk1892 n361__r_out n363__r_out 3.1
rk1894 n366__r_out n368__r_out 393.3e-3
rk1895 n368__r_out n367__r_out 5.4217
rk1896 n367__r_out n368__r_out 3.9474
rk1897 n231__vddio n232__vddio 4.884
rk1898 n232__vddio n233__vddio 1.0058
rk1899 n233__vddio n234__vddio 500.7e-3
rk1900 n234__vddio n231__vddio 4.769
rk1901 n231__vddio n232__vddio 3.1
rk1902 n231__vddio n234__vddio 3.1
rk1903 n386__vss n387__vss 4.4449
rk1904 n387__vss n386__vss 4.9153
rk1905 n369__r_out n370__r_out 4.884
rk1906 n370__r_out n371__r_out 1.5153
rk1907 n371__r_out n372__r_out 603.5e-3
rk1908 n372__r_out n369__r_out 4.1603
rk1909 n369__r_out n370__r_out 3.1
rk1910 n369__r_out n371__r_out 3.1
rk1912 n374__r_out n376__r_out 392e-3
rk1913 n376__r_out n375__r_out 5.4217
rk1914 n375__r_out n376__r_out 3.9474
rk1915 n235__vddio n236__vddio 4.884
rk1916 n236__vddio n237__vddio 1.0108
rk1917 n237__vddio n238__vddio 499.3e-3
rk1918 n238__vddio n235__vddio 4.769
rk1919 n235__vddio n236__vddio 3.1
rk1920 n235__vddio n238__vddio 3.1
rk1921 n388__vss n389__vss 4.4499
rk1922 n389__vss n388__vss 4.9139
rk1923 n377__r_out n378__r_out 4.884
rk1924 n378__r_out n379__r_out 1.5153
rk1925 n379__r_out n380__r_out 600.4e-3
rk1926 n380__r_out n377__r_out 4.1634
rk1927 n377__r_out n378__r_out 3.1
rk1928 n377__r_out n379__r_out 3.1
rk1930 n382__r_out n384__r_out 395.2e-3
rk1931 n384__r_out n383__r_out 5.4217
rk1932 n383__r_out n384__r_out 3.9474
rk1933 n239__vddio n240__vddio 4.884
rk1934 n240__vddio n241__vddio 1.0076
rk1935 n241__vddio n242__vddio 502.5e-3
rk1936 n242__vddio n239__vddio 4.769
rk1937 n239__vddio n240__vddio 3.1
rk1938 n239__vddio n242__vddio 3.1
rk1939 n390__vss n391__vss 4.4467
rk1940 n391__vss n390__vss 4.9171
rk1941 n385__r_out n386__r_out 4.884
rk1942 n386__r_out n387__r_out 1.5153
rk1943 n387__r_out n388__r_out 598.5e-3
rk1944 n388__r_out n385__r_out 4.1616
rk1945 n385__r_out n386__r_out 3.1
rk1946 n385__r_out n387__r_out 3.1
rk1948 n390__r_out n392__r_out 393.3e-3
rk1949 n392__r_out n391__r_out 5.4217
rk1950 n391__r_out n392__r_out 3.9474
rk1951 n243__vddio n244__vddio 4.884
rk1952 n244__vddio n245__vddio 1.0058
rk1953 n245__vddio n246__vddio 500.7e-3
rk1954 n246__vddio n243__vddio 4.769
rk1955 n243__vddio n244__vddio 3.1
rk1956 n243__vddio n246__vddio 3.1
rk1957 n392__vss n393__vss 4.4449
rk1958 n393__vss n392__vss 4.9153
rk1959 n393__r_out n394__r_out 4.884
rk1960 n394__r_out n395__r_out 1.5153
rk1961 n395__r_out n396__r_out 603.5e-3
rk1962 n396__r_out n393__r_out 4.1603
rk1963 n393__r_out n394__r_out 3.1
rk1964 n393__r_out n395__r_out 3.1
rk1966 n398__r_out n400__r_out 392e-3
rk1967 n400__r_out n399__r_out 5.4217
rk1968 n399__r_out n400__r_out 3.9474
rk1969 n247__vddio n248__vddio 4.884
rk1970 n248__vddio n249__vddio 1.0108
rk1971 n249__vddio n250__vddio 499.3e-3
rk1972 n250__vddio n247__vddio 4.769
rk1973 n247__vddio n248__vddio 3.1
rk1974 n247__vddio n250__vddio 3.1
rk1975 n394__vss n395__vss 4.4499
rk1976 n395__vss n394__vss 4.9139
rk1977 n361__i12__net3 n362__i12__net3 4.7406
rk1978 n362__i12__net3 n363__i12__net3 1.5153
rk1979 n363__i12__net3 n364__i12__net3 1.4995
rk1980 n364__i12__net3 n90__i12__net3 180.5e-3
rk1981 n90__i12__net3 n365__i12__net3 674.2e-3
rk1982 n365__i12__net3 n95__i12__net3 620.5e-3
rk1983 n95__i12__net3 n367__i12__net3 363.6e-3
rk1984 n367__i12__net3 n366__i12__net3 5.2385
rk1985 n365__i12__net3 n368__i12__net3 304.4e-3
rk1986 n368__i12__net3 n369__i12__net3 178.2e-3
rk1987 n369__i12__net3 n370__i12__net3 178.2e-3
rk1988 n370__i12__net3 n371__i12__net3 178.2e-3
rk1989 n371__i12__net3 n372__i12__net3 178.2e-3
rk1990 n372__i12__net3 n373__i12__net3 178.2e-3
rk1991 n373__i12__net3 n374__i12__net3 178.2e-3
rk1992 n374__i12__net3 n375__i12__net3 178.2e-3
rk1993 n375__i12__net3 n376__i12__net3 178.2e-3
rk1994 n376__i12__net3 n377__i12__net3 178.2e-3
rk1995 n377__i12__net3 n378__i12__net3 178.2e-3
rk1996 n378__i12__net3 n379__i12__net3 178.2e-3
rk1997 n379__i12__net3 n380__i12__net3 178.2e-3
rk1998 n380__i12__net3 n381__i12__net3 178.2e-3
rk1999 n381__i12__net3 n382__i12__net3 178.2e-3
rk2000 n382__i12__net3 n383__i12__net3 178.2e-3
rk2001 n383__i12__net3 n384__i12__net3 178.2e-3
rk2002 n384__i12__net3 n385__i12__net3 178.2e-3
rk2003 n385__i12__net3 n386__i12__net3 178.2e-3
rk2004 n386__i12__net3 n387__i12__net3 178.2e-3
rk2005 n387__i12__net3 n388__i12__net3 178.2e-3
rk2006 n388__i12__net3 n389__i12__net3 178.2e-3
rk2007 n389__i12__net3 n390__i12__net3 178.2e-3
rk2008 n390__i12__net3 n391__i12__net3 178.2e-3
rk2009 n391__i12__net3 n392__i12__net3 178.2e-3
rk2010 n392__i12__net3 n393__i12__net3 178.2e-3
rk2011 n393__i12__net3 n394__i12__net3 178.2e-3
rk2012 n394__i12__net3 n395__i12__net3 178.2e-3
rk2013 n395__i12__net3 n396__i12__net3 178.2e-3
rk2014 n396__i12__net3 n397__i12__net3 178.2e-3
rk2015 n397__i12__net3 n398__i12__net3 178.2e-3
rk2016 n398__i12__net3 n399__i12__net3 178.2e-3
rk2017 n399__i12__net3 n400__i12__net3 178.2e-3
rk2018 n400__i12__net3 n401__i12__net3 178.2e-3
rk2019 n401__i12__net3 n402__i12__net3 178.2e-3
rk2020 n402__i12__net3 n403__i12__net3 178.2e-3
rk2021 n403__i12__net3 n404__i12__net3 178.2e-3
rk2022 n404__i12__net3 n405__i12__net3 178.2e-3
rk2023 n405__i12__net3 n406__i12__net3 178.2e-3
rk2024 n406__i12__net3 n407__i12__net3 178.2e-3
rk2025 n407__i12__net3 n408__i12__net3 178.2e-3
rk2026 n408__i12__net3 n409__i12__net3 178.2e-3
rk2027 n409__i12__net3 n410__i12__net3 178.2e-3
rk2028 n410__i12__net3 n411__i12__net3 178.2e-3
rk2029 n411__i12__net3 n412__i12__net3 178.2e-3
rk2030 n412__i12__net3 n413__i12__net3 178.2e-3
rk2031 n413__i12__net3 n414__i12__net3 178.2e-3
rk2032 n414__i12__net3 n415__i12__net3 178.2e-3
rk2033 n415__i12__net3 n416__i12__net3 178.2e-3
rk2034 n416__i12__net3 n417__i12__net3 178.2e-3
rk2035 n417__i12__net3 n418__i12__net3 178.2e-3
rk2036 n418__i12__net3 n419__i12__net3 178.2e-3
rk2037 n419__i12__net3 n420__i12__net3 178.2e-3
rk2038 n420__i12__net3 n421__i12__net3 178.2e-3
rk2039 n421__i12__net3 n422__i12__net3 178.2e-3
rk2040 n422__i12__net3 n423__i12__net3 178.2e-3
rk2041 n423__i12__net3 n424__i12__net3 178.2e-3
rk2042 n424__i12__net3 n425__i12__net3 178.2e-3
rk2043 n425__i12__net3 n426__i12__net3 178.2e-3
rk2044 n426__i12__net3 n427__i12__net3 178.2e-3
rk2045 n427__i12__net3 n428__i12__net3 178.2e-3
rk2046 n428__i12__net3 n429__i12__net3 178.2e-3
rk2047 n429__i12__net3 n430__i12__net3 178.2e-3
rk2048 n430__i12__net3 n431__i12__net3 178.2e-3
rk2049 n431__i12__net3 n432__i12__net3 178.2e-3
rk2050 n432__i12__net3 n433__i12__net3 178.2e-3
rk2051 n433__i12__net3 n434__i12__net3 178.2e-3
rk2052 n434__i12__net3 n435__i12__net3 178.2e-3
rk2053 n435__i12__net3 n436__i12__net3 178.2e-3
rk2054 n436__i12__net3 n437__i12__net3 178.2e-3
rk2055 n437__i12__net3 n438__i12__net3 178.2e-3
rk2056 n438__i12__net3 n439__i12__net3 178.2e-3
rk2057 n439__i12__net3 n440__i12__net3 178.2e-3
rk2058 n440__i12__net3 n441__i12__net3 178.2e-3
rk2059 n441__i12__net3 n442__i12__net3 178.2e-3
rk2060 n442__i12__net3 n443__i12__net3 178.2e-3
rk2061 n443__i12__net3 n444__i12__net3 178.2e-3
rk2062 n444__i12__net3 n445__i12__net3 178.2e-3
rk2063 n445__i12__net3 n446__i12__net3 178.2e-3
rk2064 n446__i12__net3 n447__i12__net3 178.2e-3
rk2065 n447__i12__net3 n448__i12__net3 178.2e-3
rk2066 n448__i12__net3 n449__i12__net3 178.2e-3
rk2067 n449__i12__net3 n450__i12__net3 178.2e-3
rk2068 n450__i12__net3 n451__i12__net3 178.2e-3
rk2069 n451__i12__net3 n452__i12__net3 178.2e-3
rk2070 n452__i12__net3 n453__i12__net3 178.2e-3
rk2071 n453__i12__net3 n454__i12__net3 178.2e-3
rk2072 n454__i12__net3 n455__i12__net3 178.2e-3
rk2073 n455__i12__net3 n456__i12__net3 178.2e-3
rk2074 n456__i12__net3 n457__i12__net3 178.2e-3
rk2075 n457__i12__net3 n458__i12__net3 178.2e-3
rk2076 n458__i12__net3 n459__i12__net3 178.2e-3
rk2077 n459__i12__net3 n460__i12__net3 178.2e-3
rk2078 n460__i12__net3 n461__i12__net3 178.2e-3
rk2079 n461__i12__net3 n462__i12__net3 178.2e-3
rk2080 n462__i12__net3 n463__i12__net3 178.2e-3
rk2081 n463__i12__net3 n464__i12__net3 178.2e-3
rk2082 n464__i12__net3 n465__i12__net3 178.2e-3
rk2083 n465__i12__net3 n466__i12__net3 178.2e-3
rk2084 n466__i12__net3 n358__i12__net3 45.1777
rk2085 n361__i12__net3 n362__i12__net3 3.1
rk2086 n361__i12__net3 n363__i12__net3 3.1
rk2087 n361__i12__net3 n364__i12__net3 3.2632
rk2088 n366__i12__net3 n367__i12__net3 3.9474
rk2089 i12__net3 n368__i12__net3 45
rk2090 n4__i12__net3 n369__i12__net3 45
rk2091 n7__i12__net3 n370__i12__net3 45
rk2092 n20__i12__net3 n371__i12__net3 45
rk2093 n23__i12__net3 n372__i12__net3 45
rk2094 n36__i12__net3 n373__i12__net3 45
rk2095 n39__i12__net3 n374__i12__net3 45
rk2096 n52__i12__net3 n375__i12__net3 45
rk2097 n55__i12__net3 n376__i12__net3 45
rk2098 n68__i12__net3 n377__i12__net3 45
rk2099 n71__i12__net3 n378__i12__net3 45
rk2100 n84__i12__net3 n379__i12__net3 45
rk2101 n87__i12__net3 n380__i12__net3 45
rk2102 n100__i12__net3 n381__i12__net3 45
rk2103 n103__i12__net3 n382__i12__net3 45
rk2104 n106__i12__net3 n383__i12__net3 45
rk2105 n109__i12__net3 n384__i12__net3 45
rk2106 n112__i12__net3 n385__i12__net3 45
rk2107 n115__i12__net3 n386__i12__net3 45
rk2108 n118__i12__net3 n387__i12__net3 45
rk2109 n121__i12__net3 n388__i12__net3 45
rk2110 n124__i12__net3 n389__i12__net3 45
rk2111 n127__i12__net3 n390__i12__net3 45
rk2112 n130__i12__net3 n391__i12__net3 45
rk2113 n133__i12__net3 n392__i12__net3 45
rk2114 n136__i12__net3 n393__i12__net3 45
rk2115 n139__i12__net3 n394__i12__net3 45
rk2116 n142__i12__net3 n395__i12__net3 45
rk2117 n145__i12__net3 n396__i12__net3 45
rk2118 n148__i12__net3 n397__i12__net3 45
rk2119 n151__i12__net3 n398__i12__net3 45
rk2120 n154__i12__net3 n399__i12__net3 45
rk2121 n157__i12__net3 n400__i12__net3 45
rk2122 n160__i12__net3 n401__i12__net3 45
rk2123 n163__i12__net3 n402__i12__net3 45
rk2124 n166__i12__net3 n403__i12__net3 45
rk2125 n169__i12__net3 n404__i12__net3 45
rk2126 n172__i12__net3 n405__i12__net3 45
rk2127 n175__i12__net3 n406__i12__net3 45
rk2128 n178__i12__net3 n407__i12__net3 45
rk2129 n181__i12__net3 n408__i12__net3 45
rk2130 n184__i12__net3 n409__i12__net3 45
rk2131 n187__i12__net3 n410__i12__net3 45
rk2132 n190__i12__net3 n411__i12__net3 45
rk2133 n193__i12__net3 n412__i12__net3 45
rk2134 n196__i12__net3 n413__i12__net3 45
rk2135 n199__i12__net3 n414__i12__net3 45
rk2136 n202__i12__net3 n415__i12__net3 45
rk2137 n205__i12__net3 n416__i12__net3 45
rk2138 n208__i12__net3 n417__i12__net3 45
rk2139 n211__i12__net3 n418__i12__net3 45
rk2140 n214__i12__net3 n419__i12__net3 45
rk2141 n217__i12__net3 n420__i12__net3 45
rk2142 n220__i12__net3 n421__i12__net3 45
rk2143 n223__i12__net3 n422__i12__net3 45
rk2144 n226__i12__net3 n423__i12__net3 45
rk2145 n229__i12__net3 n424__i12__net3 45
rk2146 n232__i12__net3 n425__i12__net3 45
rk2147 n235__i12__net3 n426__i12__net3 45
rk2148 n238__i12__net3 n427__i12__net3 45
rk2149 n241__i12__net3 n428__i12__net3 45
rk2150 n244__i12__net3 n429__i12__net3 45
rk2151 n247__i12__net3 n430__i12__net3 45
rk2152 n250__i12__net3 n431__i12__net3 45
rk2153 n253__i12__net3 n432__i12__net3 45
rk2154 n256__i12__net3 n433__i12__net3 45
rk2155 n259__i12__net3 n434__i12__net3 45
rk2156 n262__i12__net3 n435__i12__net3 45
rk2157 n265__i12__net3 n436__i12__net3 45
rk2158 n268__i12__net3 n437__i12__net3 45
rk2159 n271__i12__net3 n438__i12__net3 45
rk2160 n274__i12__net3 n439__i12__net3 45
rk2161 n277__i12__net3 n440__i12__net3 45
rk2162 n280__i12__net3 n441__i12__net3 45
rk2163 n283__i12__net3 n442__i12__net3 45
rk2164 n286__i12__net3 n443__i12__net3 45
rk2165 n289__i12__net3 n444__i12__net3 45
rk2166 n292__i12__net3 n445__i12__net3 45
rk2167 n295__i12__net3 n446__i12__net3 45
rk2168 n298__i12__net3 n447__i12__net3 45
rk2169 n301__i12__net3 n448__i12__net3 45
rk2170 n304__i12__net3 n449__i12__net3 45
rk2171 n307__i12__net3 n450__i12__net3 45
rk2172 n310__i12__net3 n451__i12__net3 45
rk2173 n313__i12__net3 n452__i12__net3 45
rk2174 n316__i12__net3 n453__i12__net3 45
rk2175 n319__i12__net3 n454__i12__net3 45
rk2176 n322__i12__net3 n455__i12__net3 45
rk2177 n325__i12__net3 n456__i12__net3 45
rk2178 n328__i12__net3 n457__i12__net3 45
rk2179 n331__i12__net3 n458__i12__net3 45
rk2180 n334__i12__net3 n459__i12__net3 45
rk2181 n337__i12__net3 n460__i12__net3 45
rk2182 n340__i12__net3 n461__i12__net3 45
rk2183 n343__i12__net3 n462__i12__net3 45
rk2184 n346__i12__net3 n463__i12__net3 45
rk2185 n349__i12__net3 n464__i12__net3 45
rk2186 n352__i12__net3 n465__i12__net3 45
rk2187 n355__i12__net3 n466__i12__net3 45
rk2188 n7__vss n396__vss 8.0886
rk2189 n251__vddio n13__vddio 7.0956
rk2190 r_out n401__r_out 442.1e-3
rk2191 n401__r_out n402__r_out 507.8e-3
rk2192 n402__r_out n404__r_out 395.2e-3
rk2193 n404__r_out n403__r_out 5.4217
rk2194 n401__r_out n406__r_out 941.7e-3
rk2195 n406__r_out n407__r_out 900.3e-3
rk2196 n407__r_out n408__r_out 600.4e-3
rk2197 n408__r_out n409__r_out 1.5153
rk2198 n409__r_out n405__r_out 4.884
rk2199 n403__r_out n404__r_out 3.9474
rk2200 n405__r_out n406__r_out 3.2632
rk2201 n405__r_out n408__r_out 3.1
rk2202 n405__r_out n409__r_out 3.1
rl1 clkb n2__clkb 83.7904
rl2 n1__clk n2__clk 84.5404
rl3 i0__net1 n2__i0__net1 83.3077
rl4 i0__net1 n3__i0__net1 169.231
rl5 n3__clk n4__clk 56.5719
rl6 n4__clk n5__clk 48.1183
rl7 n4__clk n6__clk 56.5719
rl8 i0__net2 n2__i0__net2 82.5518
rl9 n2__i0__net2 n3__i0__net2 169.231
rl10 n3__clkb n4__clkb 83.6772
rl11 n7__clk n8__clk 88.4636
rl12 clk2 n2__clk2 112.341
rl13 n2__clk2 n3__clk2 45
rl14 n2__clk2 n4__clk2 46.9565
rl15 n5__clk2 n6__clk2 84.5404
rl16 n4__i0__net1 n5__i0__net1 84.5404
rl17 i0__net4 n2__i0__net4 86.9319
rl18 i0__net4 n3__i0__net4 169.231
rl19 i0__net6 n2__i0__net6 82.5518
rl20 n2__i0__net6 n3__i0__net6 169.231
rl21 n6__i0__net1 n7__i0__net1 83.6772
rl22 n7__clk2 n8__clk2 88.4636
rl23 i0__net3 n2__i0__net3 112.341
rl24 n2__i0__net3 n3__i0__net3 45
rl25 n2__i0__net3 n4__i0__net3 46.9565
rl26 n4__i0__net4 n5__i0__net4 112.341
rl27 n5__i0__net4 n6__i0__net4 45
rl28 n5__i0__net4 n7__i0__net4 46.9565
rl29 clk4 n2__clk4 112.341
rl30 n2__clk4 n3__clk4 45
rl31 n2__clk4 n4__clk4 46.9565
rl32 x2 n2__x2 33.7903
rl33 n2__x2 n3__x2 118.406
rl34 x0 n2__x0 33.7903
rl35 n2__x0 n3__x0 118.406
rl36 clk4b n2__clk4b 83.7904
rl37 n3__clk4b n4__clk4b 83.7904
rl38 n5__clk4 n6__clk4 84.5404
rl39 n7__clk4 n8__clk4 84.5404
rl40 y2 n2__y2 103.826
rl41 n2__y2 n3__y2 49.9799
rl42 n1__yin0 n2__yin0 85.2307
rl43 n1__yin0 n3__yin0 169.231
rl44 n1__xin0 n2__xin0 85.2307
rl45 n1__xin0 n3__xin0 169.231
rl46 y0 n2__y0 103.826
rl47 n2__y0 n3__y0 49.9799
rl48 i2__net1 n2__i2__net1 86.5999
rl49 n2__i2__net1 n3__i2__net1 169.231
rl50 i1__net1 n2__i1__net1 86.5999
rl51 n2__i1__net1 n3__i1__net1 169.231
rl52 n4__x2 n5__x2 45.0334
rl53 n5__x2 n6__x2 45
rl54 n5__x2 n7__x2 129.649
rl55 n5__clk4b n6__clk4b 83.6772
rl56 n9__clk4 n10__clk4 88.4636
rl57 n7__clk4b n8__clk4b 83.6772
rl58 n11__clk4 n12__clk4 88.4636
rl59 n4__x0 n5__x0 45.0334
rl60 n5__x0 n6__x0 45
rl61 n5__x0 n7__x0 129.649
rl62 i5__bbar n2__i5__bbar 76.9251
rl63 i5__bbar n3__i5__bbar 184.615
rl64 n1__rst n2__rst 89.4464
rl65 n3__rst n4__rst 89.4464
rl66 i3__bbar n2__i3__bbar 76.9251
rl67 i3__bbar n3__i3__bbar 184.615
rl68 i5__abar n2__i5__abar 83.3077
rl69 i5__abar n3__i5__abar 184.615
rl70 i3__abar n2__i3__abar 83.3077
rl71 i3__abar n3__i3__abar 184.615
rl72 n5__rst n6__rst 90.3096
rl73 n7__rst n8__rst 90.3096
rl74 n4__y2 n5__y2 129.649
rl75 n5__y2 n6__y2 45
rl76 n5__y2 n7__y2 45.0334
rl77 n4__y0 n5__y0 129.649
rl78 n5__y0 n6__y0 45
rl79 n5__y0 n7__y0 45.0334
rl80 i2__rstb n2__i2__rstb 79.831
rl81 i1__rstb n2__i1__rstb 79.831
rl82 n3__i2__rstb n4__i2__rstb 79.831
rl83 n3__i1__rstb n4__i1__rstb 79.831
rl84 n9__clk4b n10__clk4b 83.7904
rl85 n11__clk4b n12__clk4b 83.7904
rl86 n13__clk4 n14__clk4 84.5404
rl87 n15__clk4 n16__clk4 84.5404
rl88 n1__yin1 n2__yin1 85.2307
rl89 n1__yin1 n3__yin1 169.231
rl90 n1__xin1 n2__xin1 85.2307
rl91 n1__xin1 n3__xin1 169.231
rl92 i2__net3 n2__i2__net3 86.5999
rl93 n2__i2__net3 n3__i2__net3 169.231
rl94 i1__net3 n2__i1__net3 86.5999
rl95 n2__i1__net3 n3__i1__net3 169.231
rl96 n13__clk4b n14__clk4b 83.6772
rl97 n17__clk4 n18__clk4 88.4636
rl98 n15__clk4b n16__clk4b 83.6772
rl99 n19__clk4 n20__clk4 88.4636
rl100 n17__clk4b n18__clk4b 83.7904
rl101 n19__clk4b n20__clk4b 83.7904
rl102 n21__clk4 n22__clk4 84.5404
rl103 n23__clk4 n24__clk4 84.5404
rl104 n1__yin2 n2__yin2 85.2307
rl105 n1__yin2 n3__yin2 169.231
rl106 n1__xin2 n2__xin2 85.2307
rl107 n1__xin2 n3__xin2 169.231
rl108 i2__net4 n2__i2__net4 169.231
rl109 i2__net4 n3__i2__net4 76.6622
rl110 i1__net4 n2__i1__net4 169.231
rl111 i1__net4 n3__i1__net4 76.6622
rl112 x3 n2__x3 33.7903
rl113 n2__x3 n3__x3 118.406
rl114 n21__clk4b n22__clk4b 83.6772
rl115 n25__clk4 n26__clk4 95.2157
rl116 n23__clk4b n24__clk4b 83.6772
rl117 n27__clk4 n28__clk4 95.2157
rl118 y3 n2__y3 103.826
rl119 n2__y3 n3__y3 49.9799
rl120 n9__rst n10__rst 89.4464
rl121 n11__rst n12__rst 89.4464
rl122 n5__i2__rstb n6__i2__rstb 77.044
rl123 n5__i1__rstb n6__i1__rstb 77.044
rl124 n4__x3 n5__x3 45.0334
rl125 n5__x3 n6__x3 45
rl126 n5__x3 n7__x3 129.649
rl127 x1 n2__x1 33.7903
rl128 n2__x1 n3__x1 118.406
rl129 n25__clk4b n26__clk4b 83.7904
rl130 n27__clk4b n28__clk4b 83.7904
rl131 n29__clk4 n30__clk4 84.5404
rl132 n31__clk4 n32__clk4 84.5404
rl133 i6__bbar n2__i6__bbar 76.9251
rl134 i6__bbar n3__i6__bbar 184.615
rl135 n1__yin3 n2__yin3 85.2307
rl136 n1__yin3 n3__yin3 169.231
rl137 n1__xin3 n2__xin3 85.2307
rl138 n1__xin3 n3__xin3 169.231
rl139 y1 n2__y1 103.826
rl140 n2__y1 n3__y1 49.9799
rl141 i6__abar n2__i6__abar 83.3077
rl142 i6__abar n3__i6__abar 184.615
rl143 i2__net2 n2__i2__net2 86.5999
rl144 n2__i2__net2 n3__i2__net2 169.231
rl145 i1__net2 n2__i1__net2 86.5999
rl146 n2__i1__net2 n3__i1__net2 169.231
rl147 n4__y3 n5__y3 129.649
rl148 n5__y3 n6__y3 45
rl149 n5__y3 n7__y3 45.0334
rl150 n33__clk4b n34__clk4b 83.6772
rl151 n37__clk4 n38__clk4 88.4636
rl152 n35__clk4b n36__clk4b 83.6772
rl153 n39__clk4 n40__clk4 88.4636
rl154 n4__x1 n5__x1 45.0334
rl155 n5__x1 n6__x1 45
rl156 n5__x1 n7__x1 129.649
rl157 i4__bbar n2__i4__bbar 76.9251
rl158 i4__bbar n3__i4__bbar 184.615
rl159 n13__rst n14__rst 91.3695
rl160 n15__rst n16__rst 91.3695
rl161 i4__abar n2__i4__abar 83.3077
rl162 i4__abar n3__i4__abar 184.615
rl163 n7__i2__rstb n8__i2__rstb 79.9443
rl164 n7__i1__rstb n8__i1__rstb 79.9443
rl165 n21__rst n22__rst 110.418
rl166 n22__rst n23__rst 45
rl167 n22__rst n24__rst 48.8796
rl168 n25__rst n26__rst 110.418
rl169 n26__rst n27__rst 45
rl170 n26__rst n28__rst 48.8796
rl171 n7__y1 n8__y1 129.649
rl172 n8__y1 n9__y1 45
rl173 n8__y1 n10__y1 45.0334
rl174 n5__a2 n6__a2 53.079
rl175 n6__a2 n7__a2 87.6944
rl176 n7__a2 n8__a2 144.231
rl177 n8__a2 n9__a2 94.2308
rl178 n5__a0 n6__a0 53.079
rl179 n6__a0 n7__a0 87.6944
rl180 n7__a0 n8__a0 144.231
rl181 n8__a0 n9__a0 94.2308
rl182 a3 n2__a3 108.848
rl183 n2__a3 n3__a3 31.9251
rl184 n3__a3 n4__a3 144.231
rl185 n4__a3 n5__a3 94.2308
rl186 a1 n2__a1 108.848
rl187 n2__a1 n3__a1 31.9251
rl188 n3__a1 n4__a1 144.231
rl189 n4__a1 n5__a1 94.2308
rl190 i8__net51 n2__i8__net51 205.002
rl191 n2__i8__net51 n3__i8__net51 264.617
rl192 i7__net51 n2__i7__net51 205.002
rl193 n2__i7__net51 n3__i7__net51 264.617
rl194 i8__carry_bar n2__i8__carry_bar 181.925
rl195 n2__i8__carry_bar n3__i8__carry_bar 380.002
rl196 i7__carry_bar n2__i7__carry_bar 181.925
rl197 n2__i7__carry_bar n3__i7__carry_bar 380.002
rl198 n10__a2 n11__a2 85.7713
rl199 n11__a2 n12__a2 476.156
rl200 n10__a0 n11__a0 85.7713
rl201 n11__a0 n12__a0 476.156
rl202 n6__a3 n7__a3 205.223
rl203 n7__a3 n8__a3 360.993
rl204 n6__a1 n7__a1 205.223
rl205 n7__a1 n8__a1 360.993
rl206 c0 n2__c0 91.1873
rl207 n2__c0 n3__c0 48.1183
rl208 n2__c0 n4__c0 229.649
rl209 c1 n2__c1 137.341
rl210 n2__c1 n3__c1 47.4801
rl211 n2__c1 n4__c1 183.495
rl212 s0 n2__s0 53.079
rl213 n2__s0 n3__s0 87.6944
rl214 n3__s0 n4__s0 144.231
rl215 n4__s0 n5__s0 94.2308
rl216 net12 n2__net12 198.88
rl217 n2__net12 n3__net12 46.8551
rl218 n2__net12 n4__net12 102.726
rl219 s1 n2__s1 108.848
rl220 n2__s1 n3__s1 31.9251
rl221 n3__s1 n4__s1 144.231
rl222 n4__s1 n5__s1 94.2308
rl223 n5__c0 n6__c0 83.495
rl224 n6__c0 n7__c0 47.4801
rl225 n6__c0 n8__c0 218.11
rl226 n5__c1 n6__c1 129.649
rl227 n6__c1 n7__c1 48.1183
rl228 n6__c1 n8__c1 171.957
rl229 i9__net51 n2__i9__net51 205.002
rl230 n2__i9__net51 n3__i9__net51 264.617
rl231 i10__net116 n2__i10__net116 260.418
rl232 n2__i10__net116 n3__i10__net116 48.1183
rl233 n2__i10__net116 n4__i10__net116 41.1873
rl234 i9__carry_bar n2__i9__carry_bar 181.925
rl235 n2__i9__carry_bar n3__i9__carry_bar 380.002
rl236 n5__net12 n6__net12 202.726
rl237 n6__net12 n7__net12 47.4801
rl238 n6__net12 n8__net12 98.8796
rl239 n9__c1 n10__c1 129.649
rl240 n10__c1 n11__c1 46.8551
rl241 n10__c1 n12__c1 171.957
rl242 n6__s0 n7__s0 85.7713
rl243 n7__s0 n8__s0 476.156
rl244 n9__c0 n10__c0 83.495
rl245 n10__c0 n11__c0 47.4801
rl246 n10__c0 n12__c0 218.11
rl247 n6__s1 n7__s1 205.223
rl248 n7__s1 n8__s1 360.993
rl249 n9__net12 n10__net12 202.726
rl250 n10__net12 n11__net12 48.1183
rl251 n10__net12 n12__net12 98.8796
rl252 n13__c1 n14__c1 152.726
rl253 n14__c1 n15__c1 47.4801
rl254 n14__c1 n16__c1 148.88
rl255 n13__c0 n14__c0 83.495
rl256 n14__c0 n15__c0 46.8551
rl257 n14__c0 n16__c0 218.11
rl258 i10__net114 n2__i10__net114 147.465
rl259 n2__i10__net114 n3__i10__net114 311.538
rl260 n3__i10__net114 n4__i10__net114 45.0334
rl262 n4__i10__net114 n6__i10__net114 47.4801
rl263 n5__i10__net116 n6__i10__net116 260.418
rl264 n6__i10__net116 n7__i10__net116 45
rl265 n6__i10__net116 n8__i10__net116 41.1873
rl266 n69__clk4 n70__clk4 85.3076
rl267 n70__clk4 n71__clk4 62.2307
rl268 n17__clk2 n18__clk2 85.9926
rl269 n18__clk2 n19__clk2 62.9157
rl270 n45__rst n46__rst 45
rl271 n46__rst n47__rst 48.8796
rl272 n46__rst n48__rst 110.418
rl273 i14__i3__rstb n2__i14__i3__rstb 79.081
rl274 i14__i7__net1 n2__i14__i7__net1 90.0987
rl275 n2__i14__i7__net1 n3__i14__i7__net1 45.5166
rl276 n2__i14__i7__net1 n4__i14__i7__net1 74.7141
rl277 n49__rst n50__rst 92.2327
rl278 n15__clk n16__clk 88.4636
rl279 n12__clkb n13__clkb 84.5404
rl280 i14__i3__net5 n2__i14__i3__net5 75.2349
rl281 i14__i3__net5 n3__i14__i3__net5 169.231
rl282 i14__net2 n2__i14__net2 85.2307
rl283 n2__i14__net2 n3__i14__net2 169.231
rl284 n17__clk n18__clk 83.6772
rl285 n14__clkb n15__clkb 82.9272
rl286 i14__shift n2__i14__shift 124.714
rl287 n2__i14__shift n3__i14__shift 50.1123
rl288 n2__i14__shift n4__i14__shift 40.0987
rl289 n51__rst n52__rst 45
rl290 n52__rst n53__rst 48.8796
rl291 n52__rst n54__rst 110.418
rl292 i14__i4__rstb n2__i14__i4__rstb 79.081
rl293 i14__i0__net1 n2__i14__i0__net1 88.6964
rl294 n5__i14__shift n6__i14__shift 86.0764
rl295 n55__rst n56__rst 92.2327
rl296 n3__i14__i0__net1 n4__i14__i0__net1 69.5191
rl297 n7__i14__shift n8__i14__shift 114.773
rl298 n19__clk n20__clk 88.4636
rl299 n16__clkb n17__clkb 84.5404
rl300 i14__i4__net5 n2__i14__i4__net5 75.2349
rl301 i14__i4__net5 n3__i14__i4__net5 169.231
rl302 n9__i14__shift n10__i14__shift 124.714
rl303 n10__i14__shift n11__i14__shift 50.1123
rl304 n10__i14__shift n12__i14__shift 40.0987
rl305 i14__net8 n2__i14__net8 85.2307
rl306 n2__i14__net8 n3__i14__net8 169.231
rl307 n21__clk n22__clk 83.6772
rl308 n18__clkb n19__clkb 82.9272
rl309 i14__i1__net1 n2__i14__i1__net1 88.6964
rl310 n13__i14__shift n14__i14__shift 86.0764
rl311 n3__i14__i1__net1 n4__i14__i1__net1 69.5191
rl312 n15__i14__shift n16__i14__shift 114.773
rl313 n57__rst n58__rst 45
rl314 n58__rst n59__rst 48.8796
rl315 n58__rst n60__rst 110.418
rl316 i14__i5__rstb n2__i14__i5__rstb 79.081
rl317 n61__rst n62__rst 92.2327
rl318 n17__i14__shift n18__i14__shift 124.714
rl319 n18__i14__shift n19__i14__shift 50.1123
rl320 n18__i14__shift n20__i14__shift 40.0987
rl321 n23__clk n24__clk 88.4636
rl322 n20__clkb n21__clkb 84.5404
rl323 i14__i2__net1 n2__i14__i2__net1 88.6964
rl324 n21__i14__shift n22__i14__shift 86.0764
rl325 i14__i5__net5 n2__i14__i5__net5 75.2349
rl326 i14__i5__net5 n3__i14__i5__net5 169.231
rl327 n3__i14__i2__net1 n4__i14__i2__net1 69.5191
rl328 n23__i14__shift n24__i14__shift 114.773
rl329 i14__net14 n2__i14__net14 85.2307
rl330 n2__i14__net14 n3__i14__net14 169.231
rl331 n25__clk n26__clk 83.6772
rl332 n22__clkb n23__clkb 82.9272
rl333 r_in n2__r_in 67.0474
rl334 serial_out n2__serial_out 83.1933
rl335 net5 n2__net5 81.1099
rl336 i11__net1 n2__i11__net1 62.713
rl337 n3__serial_out n4__serial_out 116.37
rl338 n3__serial_out n5__serial_out 111.538
rl339 n3__r_in n4__r_in 29.9319
rl340 n3__r_in n5__r_in 25.7653
rl341 i12__net1 n2__i12__net1 40.3486
rl342 i12__net1 n3__i12__net1 15.3486
rl343 n4__i12__net1 n5__i12__net1 40.3486
rl344 n4__i12__net1 n6__i12__net1 15.3486
rl345 i12__net2 n2__i12__net2 40.3486
rl346 i12__net2 n3__i12__net2 15.3486
rl347 n4__i12__net2 n5__i12__net2 40.3486
rl348 n4__i12__net2 n6__i12__net2 15.3486
rl349 n7__i12__net2 n8__i12__net2 40.3486
rl350 n7__i12__net2 n9__i12__net2 15.3486
rl351 n10__i12__net2 n11__i12__net2 40.3486
rl352 n10__i12__net2 n12__i12__net2 15.3486
rl353 n13__i12__net2 n14__i12__net2 40.3486
rl354 n13__i12__net2 n15__i12__net2 15.3486
rl355 n16__i12__net2 n17__i12__net2 40.3486
rl356 n16__i12__net2 n18__i12__net2 15.3486
rl357 n19__i12__net2 n20__i12__net2 40.3486
rl358 n19__i12__net2 n21__i12__net2 15.3486
rl359 n22__i12__net2 n23__i12__net2 40.3486
rl360 n22__i12__net2 n24__i12__net2 15.3486
rl361 n25__i12__net2 n26__i12__net2 40.3486
rl362 n25__i12__net2 n27__i12__net2 15.3486
rl363 n28__i12__net2 n29__i12__net2 40.3486
rl364 n28__i12__net2 n30__i12__net2 15.3486
rl365 n38__i12__net2 n39__i12__net2 40.3486
rl366 n38__i12__net2 n40__i12__net2 15.3486
rl367 i12__net3 n2__i12__net3 40.3486
rl368 i12__net3 n3__i12__net3 15.3486
rl369 n4__i12__net3 n5__i12__net3 40.3486
rl370 n4__i12__net3 n6__i12__net3 15.3486
rl371 n7__i12__net3 n8__i12__net3 40.3486
rl372 n7__i12__net3 n9__i12__net3 15.3486
rl373 n20__i12__net3 n21__i12__net3 40.3486
rl374 n20__i12__net3 n22__i12__net3 15.3486
rl375 n23__i12__net3 n24__i12__net3 40.3486
rl376 n23__i12__net3 n25__i12__net3 15.3486
rl377 n36__i12__net3 n37__i12__net3 40.3486
rl378 n36__i12__net3 n38__i12__net3 15.3486
rl379 n39__i12__net3 n40__i12__net3 40.3486
rl380 n39__i12__net3 n41__i12__net3 15.3486
rl381 n52__i12__net3 n53__i12__net3 40.3486
rl382 n52__i12__net3 n54__i12__net3 15.3486
rl383 n55__i12__net3 n56__i12__net3 40.3486
rl384 n55__i12__net3 n57__i12__net3 15.3486
rl385 n68__i12__net3 n69__i12__net3 40.3486
rl386 n68__i12__net3 n70__i12__net3 15.3486
rl387 n71__i12__net3 n72__i12__net3 40.3486
rl388 n71__i12__net3 n73__i12__net3 15.3486
rl389 n84__i12__net3 n85__i12__net3 40.3486
rl390 n84__i12__net3 n86__i12__net3 15.3486
rl391 n87__i12__net3 n88__i12__net3 40.3486
rl392 n87__i12__net3 n89__i12__net3 15.3486
rl393 n100__i12__net3 n101__i12__net3 40.3486
rl394 n100__i12__net3 n102__i12__net3 15.3486
rl395 n103__i12__net3 n104__i12__net3 40.3486
rl396 n103__i12__net3 n105__i12__net3 15.3486
rl397 n106__i12__net3 n107__i12__net3 40.3486
rl398 n106__i12__net3 n108__i12__net3 15.3486
rl399 n109__i12__net3 n110__i12__net3 40.3486
rl400 n109__i12__net3 n111__i12__net3 15.3486
rl401 n112__i12__net3 n113__i12__net3 40.3486
rl402 n112__i12__net3 n114__i12__net3 15.3486
rl403 n115__i12__net3 n116__i12__net3 40.3486
rl404 n115__i12__net3 n117__i12__net3 15.3486
rl405 n118__i12__net3 n119__i12__net3 40.3486
rl406 n118__i12__net3 n120__i12__net3 15.3486
rl407 n121__i12__net3 n122__i12__net3 40.3486
rl408 n121__i12__net3 n123__i12__net3 15.3486
rl409 n124__i12__net3 n125__i12__net3 40.3486
rl410 n124__i12__net3 n126__i12__net3 15.3486
rl411 n127__i12__net3 n128__i12__net3 40.3486
rl412 n127__i12__net3 n129__i12__net3 15.3486
rl413 n130__i12__net3 n131__i12__net3 40.3486
rl414 n130__i12__net3 n132__i12__net3 15.3486
rl415 n133__i12__net3 n134__i12__net3 40.3486
rl416 n133__i12__net3 n135__i12__net3 15.3486
rl417 n136__i12__net3 n137__i12__net3 40.3486
rl418 n136__i12__net3 n138__i12__net3 15.3486
rl419 n139__i12__net3 n140__i12__net3 40.3486
rl420 n139__i12__net3 n141__i12__net3 15.3486
rl421 n142__i12__net3 n143__i12__net3 40.3486
rl422 n142__i12__net3 n144__i12__net3 15.3486
rl423 n145__i12__net3 n146__i12__net3 40.3486
rl424 n145__i12__net3 n147__i12__net3 15.3486
rl425 n148__i12__net3 n149__i12__net3 40.3486
rl426 n148__i12__net3 n150__i12__net3 15.3486
rl427 n151__i12__net3 n152__i12__net3 40.3486
rl428 n151__i12__net3 n153__i12__net3 15.3486
rl429 n154__i12__net3 n155__i12__net3 40.3486
rl430 n154__i12__net3 n156__i12__net3 15.3486
rl431 n157__i12__net3 n158__i12__net3 40.3486
rl432 n157__i12__net3 n159__i12__net3 15.3486
rl433 n160__i12__net3 n161__i12__net3 40.3486
rl434 n160__i12__net3 n162__i12__net3 15.3486
rl435 n163__i12__net3 n164__i12__net3 40.3486
rl436 n163__i12__net3 n165__i12__net3 15.3486
rl437 n166__i12__net3 n167__i12__net3 40.3486
rl438 n166__i12__net3 n168__i12__net3 15.3486
rl439 n169__i12__net3 n170__i12__net3 40.3486
rl440 n169__i12__net3 n171__i12__net3 15.3486
rl441 n172__i12__net3 n173__i12__net3 40.3486
rl442 n172__i12__net3 n174__i12__net3 15.3486
rl443 n175__i12__net3 n176__i12__net3 40.3486
rl444 n175__i12__net3 n177__i12__net3 15.3486
rl445 n178__i12__net3 n179__i12__net3 40.3486
rl446 n178__i12__net3 n180__i12__net3 15.3486
rl447 n181__i12__net3 n182__i12__net3 40.3486
rl448 n181__i12__net3 n183__i12__net3 15.3486
rl449 n184__i12__net3 n185__i12__net3 40.3486
rl450 n184__i12__net3 n186__i12__net3 15.3486
rl451 n187__i12__net3 n188__i12__net3 40.3486
rl452 n187__i12__net3 n189__i12__net3 15.3486
rl453 n190__i12__net3 n191__i12__net3 40.3486
rl454 n190__i12__net3 n192__i12__net3 15.3486
rl455 n193__i12__net3 n194__i12__net3 40.3486
rl456 n193__i12__net3 n195__i12__net3 15.3486
rl457 n196__i12__net3 n197__i12__net3 40.3486
rl458 n196__i12__net3 n198__i12__net3 15.3486
rl459 n199__i12__net3 n200__i12__net3 40.3486
rl460 n199__i12__net3 n201__i12__net3 15.3486
rl461 n202__i12__net3 n203__i12__net3 40.3486
rl462 n202__i12__net3 n204__i12__net3 15.3486
rl463 n205__i12__net3 n206__i12__net3 40.3486
rl464 n205__i12__net3 n207__i12__net3 15.3486
rl465 n208__i12__net3 n209__i12__net3 40.3486
rl466 n208__i12__net3 n210__i12__net3 15.3486
rl467 n211__i12__net3 n212__i12__net3 40.3486
rl468 n211__i12__net3 n213__i12__net3 15.3486
rl469 n214__i12__net3 n215__i12__net3 40.3486
rl470 n214__i12__net3 n216__i12__net3 15.3486
rl471 n217__i12__net3 n218__i12__net3 40.3486
rl472 n217__i12__net3 n219__i12__net3 15.3486
rl473 n220__i12__net3 n221__i12__net3 40.3486
rl474 n220__i12__net3 n222__i12__net3 15.3486
rl475 n223__i12__net3 n224__i12__net3 40.3486
rl476 n223__i12__net3 n225__i12__net3 15.3486
rl477 n226__i12__net3 n227__i12__net3 40.3486
rl478 n226__i12__net3 n228__i12__net3 15.3486
rl479 n229__i12__net3 n230__i12__net3 40.3486
rl480 n229__i12__net3 n231__i12__net3 15.3486
rl481 n232__i12__net3 n233__i12__net3 40.3486
rl482 n232__i12__net3 n234__i12__net3 15.3486
rl483 n235__i12__net3 n236__i12__net3 40.3486
rl484 n235__i12__net3 n237__i12__net3 15.3486
rl485 n238__i12__net3 n239__i12__net3 40.3486
rl486 n238__i12__net3 n240__i12__net3 15.3486
rl487 n241__i12__net3 n242__i12__net3 40.3486
rl488 n241__i12__net3 n243__i12__net3 15.3486
rl489 n244__i12__net3 n245__i12__net3 40.3486
rl490 n244__i12__net3 n246__i12__net3 15.3486
rl491 n247__i12__net3 n248__i12__net3 40.3486
rl492 n247__i12__net3 n249__i12__net3 15.3486
rl493 n250__i12__net3 n251__i12__net3 40.3486
rl494 n250__i12__net3 n252__i12__net3 15.3486
rl495 n253__i12__net3 n254__i12__net3 40.3486
rl496 n253__i12__net3 n255__i12__net3 15.3486
rl497 n256__i12__net3 n257__i12__net3 40.3486
rl498 n256__i12__net3 n258__i12__net3 15.3486
rl499 n259__i12__net3 n260__i12__net3 40.3486
rl500 n259__i12__net3 n261__i12__net3 15.3486
rl501 n262__i12__net3 n263__i12__net3 40.3486
rl502 n262__i12__net3 n264__i12__net3 15.3486
rl503 n265__i12__net3 n266__i12__net3 40.3486
rl504 n265__i12__net3 n267__i12__net3 15.3486
rl505 n268__i12__net3 n269__i12__net3 40.3486
rl506 n268__i12__net3 n270__i12__net3 15.3486
rl507 n271__i12__net3 n272__i12__net3 40.3486
rl508 n271__i12__net3 n273__i12__net3 15.3486
rl509 n274__i12__net3 n275__i12__net3 40.3486
rl510 n274__i12__net3 n276__i12__net3 15.3486
rl511 n277__i12__net3 n278__i12__net3 40.3486
rl512 n277__i12__net3 n279__i12__net3 15.3486
rl513 n280__i12__net3 n281__i12__net3 40.3486
rl514 n280__i12__net3 n282__i12__net3 15.3486
rl515 n283__i12__net3 n284__i12__net3 40.3486
rl516 n283__i12__net3 n285__i12__net3 15.3486
rl517 n286__i12__net3 n287__i12__net3 40.3486
rl518 n286__i12__net3 n288__i12__net3 15.3486
rl519 n289__i12__net3 n290__i12__net3 40.3486
rl520 n289__i12__net3 n291__i12__net3 15.3486
rl521 n292__i12__net3 n293__i12__net3 40.3486
rl522 n292__i12__net3 n294__i12__net3 15.3486
rl523 n295__i12__net3 n296__i12__net3 40.3486
rl524 n295__i12__net3 n297__i12__net3 15.3486
rl525 n298__i12__net3 n299__i12__net3 40.3486
rl526 n298__i12__net3 n300__i12__net3 15.3486
rl527 n301__i12__net3 n302__i12__net3 40.3486
rl528 n301__i12__net3 n303__i12__net3 15.3486
rl529 n304__i12__net3 n305__i12__net3 40.3486
rl530 n304__i12__net3 n306__i12__net3 15.3486
rl531 n307__i12__net3 n308__i12__net3 40.3486
rl532 n307__i12__net3 n309__i12__net3 15.3486
rl533 n310__i12__net3 n311__i12__net3 40.3486
rl534 n310__i12__net3 n312__i12__net3 15.3486
rl535 n313__i12__net3 n314__i12__net3 40.3486
rl536 n313__i12__net3 n315__i12__net3 15.3486
rl537 n316__i12__net3 n317__i12__net3 40.3486
rl538 n316__i12__net3 n318__i12__net3 15.3486
rl539 n319__i12__net3 n320__i12__net3 40.3486
rl540 n319__i12__net3 n321__i12__net3 15.3486
rl541 n322__i12__net3 n323__i12__net3 40.3486
rl542 n322__i12__net3 n324__i12__net3 15.3486
rl543 n325__i12__net3 n326__i12__net3 40.3486
rl544 n325__i12__net3 n327__i12__net3 15.3486
rl545 n328__i12__net3 n329__i12__net3 40.3486
rl546 n328__i12__net3 n330__i12__net3 15.3486
rl547 n331__i12__net3 n332__i12__net3 40.3486
rl548 n331__i12__net3 n333__i12__net3 15.3486
rl549 n334__i12__net3 n335__i12__net3 40.3486
rl550 n334__i12__net3 n336__i12__net3 15.3486
rl551 n337__i12__net3 n338__i12__net3 40.3486
rl552 n337__i12__net3 n339__i12__net3 15.3486
rl553 n340__i12__net3 n341__i12__net3 40.3486
rl554 n340__i12__net3 n342__i12__net3 15.3486
rl555 n343__i12__net3 n344__i12__net3 40.3486
rl556 n343__i12__net3 n345__i12__net3 15.3486
rl557 n346__i12__net3 n347__i12__net3 40.3486
rl558 n346__i12__net3 n348__i12__net3 15.3486
rl559 n349__i12__net3 n350__i12__net3 40.3486
rl560 n349__i12__net3 n351__i12__net3 15.3486
rl561 n352__i12__net3 n353__i12__net3 40.3486
rl562 n352__i12__net3 n354__i12__net3 15.3486
rl563 n355__i12__net3 n356__i12__net3 40.3486
rl564 n355__i12__net3 n357__i12__net3 15.3486
rl565 n358__i12__net3 n359__i12__net3 40.3486
rl566 n358__i12__net3 n360__i12__net3 15.3486
mi12__m5_99__rcx n239__vddio n345__i12__net3 n377__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_98__rcx n385__r_out n348__i12__net3 n239__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_97__rcx n243__vddio n351__i12__net3 n385__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_96__rcx n393__r_out n354__i12__net3 n243__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_95__rcx n247__vddio n357__i12__net3 n393__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_94__rcx n405__r_out n360__i12__net3 n247__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.3995e-12 AS=1.3995e-12 PD=19.01e-6 PS=19.01e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_93__rcx n227__vddio n327__i12__net3 n353__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_92__rcx n361__r_out n330__i12__net3 n227__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_91__rcx n231__vddio n333__i12__net3 n361__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_90__rcx n369__r_out n336__i12__net3 n231__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_89__rcx n235__vddio n339__i12__net3 n369__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_88__rcx n377__r_out n342__i12__net3 n235__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_87__rcx n353__r_out n324__i12__net3 n223__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_86__rcx n329__r_out n306__i12__net3 n211__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_85__rcx n215__vddio n309__i12__net3 n329__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_84__rcx n337__r_out n312__i12__net3 n215__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_83__rcx n219__vddio n315__i12__net3 n337__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_82__rcx n345__r_out n318__i12__net3 n219__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_81__rcx n223__vddio n321__i12__net3 n345__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_80__rcx n305__r_out n288__i12__net3 n199__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_79__rcx n203__vddio n291__i12__net3 n305__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_78__rcx n313__r_out n294__i12__net3 n203__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_77__rcx n207__vddio n297__i12__net3 n313__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_76__rcx n321__r_out n300__i12__net3 n207__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_75__rcx n211__vddio n303__i12__net3 n321__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_74__rcx n281__r_out n270__i12__net3 n187__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_73__rcx n191__vddio n273__i12__net3 n281__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_72__rcx n289__r_out n276__i12__net3 n191__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_71__rcx n195__vddio n279__i12__net3 n289__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_70__rcx n297__r_out n282__i12__net3 n195__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_69__rcx n199__vddio n285__i12__net3 n297__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_68__rcx n257__r_out n252__i12__net3 n175__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_67__rcx n179__vddio n255__i12__net3 n257__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_66__rcx n265__r_out n258__i12__net3 n179__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_65__rcx n183__vddio n261__i12__net3 n265__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_64__rcx n273__r_out n264__i12__net3 n183__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_63__rcx n187__vddio n267__i12__net3 n273__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_62__rcx n175__vddio n249__i12__net3 n249__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_61__rcx n163__vddio n231__i12__net3 n225__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_60__rcx n233__r_out n234__i12__net3 n163__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_59__rcx n167__vddio n237__i12__net3 n233__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_58__rcx n241__r_out n240__i12__net3 n167__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_57__rcx n171__vddio n243__i12__net3 n241__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_56__rcx n249__r_out n246__i12__net3 n171__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_55__rcx n151__vddio n213__i12__net3 n201__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_54__rcx n209__r_out n216__i12__net3 n151__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_53__rcx n155__vddio n219__i12__net3 n209__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_52__rcx n217__r_out n222__i12__net3 n155__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_51__rcx n159__vddio n225__i12__net3 n217__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_50__rcx n225__r_out n228__i12__net3 n159__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_49__rcx n139__vddio n195__i12__net3 n181__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_48__rcx n185__r_out n198__i12__net3 n139__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_47__rcx n143__vddio n201__i12__net3 n185__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_46__rcx n193__r_out n204__i12__net3 n143__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_45__rcx n147__vddio n207__i12__net3 n193__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_44__rcx n201__r_out n210__i12__net3 n147__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_43__rcx n126__vddio n177__i12__net3 n153__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_42__rcx n161__r_out n180__i12__net3 n126__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_41__rcx n130__vddio n183__i12__net3 n161__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_40__rcx n169__r_out n186__i12__net3 n130__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_39__rcx n134__vddio n189__i12__net3 n169__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_38__rcx n181__r_out n192__i12__net3 n134__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_37__rcx n153__r_out n174__i12__net3 n122__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_36__rcx n129__r_out n156__i12__net3 n110__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_35__rcx n114__vddio n159__i12__net3 n129__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_34__rcx n137__r_out n162__i12__net3 n114__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_33__rcx n118__vddio n165__i12__net3 n137__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_32__rcx n145__r_out n168__i12__net3 n118__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_31__rcx n122__vddio n171__i12__net3 n145__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_30__rcx n105__r_out n138__i12__net3 n98__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_29__rcx n102__vddio n141__i12__net3 n105__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_28__rcx n113__r_out n144__i12__net3 n102__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_27__rcx n106__vddio n147__i12__net3 n113__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_26__rcx n121__r_out n150__i12__net3 n106__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_25__rcx n110__vddio n153__i12__net3 n121__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_24__rcx n81__r_out n120__i12__net3 n86__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_23__rcx n90__vddio n123__i12__net3 n81__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_22__rcx n89__r_out n126__i12__net3 n90__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_21__rcx n94__vddio n129__i12__net3 n89__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_20__rcx n97__r_out n132__i12__net3 n94__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_19__rcx n98__vddio n135__i12__net3 n97__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_18__rcx n57__r_out n102__i12__net3 n74__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_17__rcx n78__vddio n105__i12__net3 n57__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_16__rcx n65__r_out n108__i12__net3 n78__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_15__rcx n82__vddio n111__i12__net3 n65__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_14__rcx n73__r_out n114__i12__net3 n82__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_13__rcx n86__vddio n117__i12__net3 n73__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_12__rcx n74__vddio n89__i12__net3 n49__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_11__rcx n62__vddio n41__i12__net3 n25__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_10__rcx n33__r_out n54__i12__net3 n62__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_9__rcx n66__vddio n57__i12__net3 n33__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_8__rcx n41__r_out n70__i12__net3 n66__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_7__rcx n70__vddio n73__i12__net3 n41__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_6__rcx n49__r_out n86__i12__net3 n70__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_5__rcx n9__r_out n6__i12__net3 n50__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_4__rcx n54__vddio n9__i12__net3 n9__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_3__rcx n17__r_out n22__i12__net3 n54__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_2__rcx n58__vddio n25__i12__net3 n17__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5_1__rcx n25__r_out n38__i12__net3 n58__vddio n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.06e-6 PS=19.06e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m5 n50__vddio n3__i12__net3 n1__r_out n13__vddio g45p2svt L=150e-9 W=9.33e-6 AD=1.866e-12 AS=1.866e-12 PD=19.01e-6 PS=19.01e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m2_10__rcx n42__i12__net3 n15__i12__net2 n30__vddio n13__vddio g45p2svt L=150e-9 W=9.43e-6 AD=1.886e-12 AS=1.886e-12 PD=19.26e-6 PS=19.26e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m2_9__rcx n34__vddio n18__i12__net2 n42__i12__net3 n13__vddio g45p2svt L=150e-9 W=9.43e-6 AD=1.886e-12 AS=1.886e-12 PD=19.26e-6 PS=19.26e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m2_8__rcx n58__i12__net3 n21__i12__net2 n34__vddio n13__vddio g45p2svt L=150e-9 W=9.43e-6 AD=1.886e-12 AS=1.886e-12 PD=19.26e-6 PS=19.26e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m2_7__rcx n38__vddio n24__i12__net2 n58__i12__net3 n13__vddio g45p2svt L=150e-9 W=9.43e-6 AD=1.886e-12 AS=1.886e-12 PD=19.26e-6 PS=19.26e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m2_6__rcx n74__i12__net3 n27__i12__net2 n38__vddio n13__vddio g45p2svt L=150e-9 W=9.43e-6 AD=1.886e-12 AS=1.886e-12 PD=19.26e-6 PS=19.26e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m2_5__rcx n42__vddio n30__i12__net2 n74__i12__net3 n13__vddio g45p2svt L=150e-9 W=9.43e-6 AD=1.886e-12 AS=1.886e-12 PD=19.26e-6 PS=19.26e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m2_4__rcx n361__i12__net3 n40__i12__net2 n42__vddio n13__vddio g45p2svt L=150e-9 W=9.43e-6 AD=1.4145e-12 AS=1.4145e-12 PD=19.21e-6 PS=19.21e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi11__m6 n2__vddio n2__r_in n5__net5 n4__vddio g45p2svt L=150e-9 W=640e-9 AD=128e-15 AS=128e-15 PD=1.63e-6 PS=1.63e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi11__m2 n6__r_in n2__net5 n2__vddio n4__vddio g45p2svt L=150e-9 W=640e-9 AD=96e-15 AS=96e-15 PD=1.63e-6 PS=1.63e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m6 n7__i12__net1 n5__r_in n25__vddio n13__vddio g45p2svt L=150e-9 W=1.28e-6 AD=192e-15 AS=192e-15 PD=2.86e-6 PS=2.86e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m1_1__rcx n21__vddio n3__i12__net1 n31__i12__net2 n13__vddio g45p2svt L=150e-9 W=5.76e-6 AD=1.152e-12 AS=1.152e-12 PD=11.87e-6 PS=11.87e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m1 n43__i12__net2 n6__i12__net1 n21__vddio n13__vddio g45p2svt L=150e-9 W=5.76e-6 AD=864e-15 AS=864e-15 PD=11.87e-6 PS=11.87e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m2_3__rcx n10__i12__net3 n3__i12__net2 n15__vddio n13__vddio g45p2svt L=150e-9 W=9.43e-6 AD=1.886e-12 AS=1.886e-12 PD=19.21e-6 PS=19.21e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m2_2__rcx n26__vddio n6__i12__net2 n10__i12__net3 n13__vddio g45p2svt L=150e-9 W=9.43e-6 AD=1.886e-12 AS=1.886e-12 PD=19.26e-6 PS=19.26e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m2_1__rcx n26__i12__net3 n9__i12__net2 n26__vddio n13__vddio g45p2svt L=150e-9 W=9.43e-6 AD=1.886e-12 AS=1.886e-12 PD=19.26e-6 PS=19.26e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m2 n30__vddio n12__i12__net2 n26__i12__net3 n13__vddio g45p2svt L=150e-9 W=9.43e-6 AD=1.886e-12 AS=1.886e-12 PD=19.26e-6 PS=19.26e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi6__pm0 n61__vdd x3 n4__i6__abar n76__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi6__pm1 n4__i6__bbar y3 n61__vdd n76__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi6__pm2 i6__net1 n4__x3 n63__vdd n76__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi6__pm3 n12__a3 i6__bbar i6__net1 n76__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi6__pm5 i6__net2 i6__abar n12__a3 n76__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi6__pm4 n74__vdd n4__y3 i6__net2 n76__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__pm0 n14__vdd x2 n4__i5__abar n57__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__pm1 n4__i5__bbar y2 n14__vdd n57__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__pm2 i5__net1 n4__x2 n18__vdd n57__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__pm3 a2 i5__bbar i5__net1 n57__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__pm5 i5__net2 i5__abar a2 n57__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__pm4 n55__vdd n4__y2 i5__net2 n57__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi4__pm0 n70__vdd x1 n4__i4__abar n139__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi4__pm1 n4__i4__bbar y1 n70__vdd n139__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi4__pm2 i4__net1 n4__x1 n72__vdd n139__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi4__pm3 n9__a1 i4__bbar i4__net1 n139__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi4__pm5 i4__net2 i4__abar n9__a1 n139__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi4__pm4 n138__vdd n7__y1 i4__net2 n139__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi3__pm0 n16__vdd x0 n4__i3__abar n60__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi3__pm1 n4__i3__bbar y0 n16__vdd n60__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi3__pm2 i3__net1 n4__x0 n20__vdd n60__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi3__pm3 a0 i3__bbar i3__net1 n60__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi3__pm5 i3__net2 i3__abar a0 n60__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi3__pm4 n58__vdd n4__y0 i3__net2 n60__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi15__pm0 n9__clkb n3__clk n5__vdd n7__vdd g45p1svt L=45e-9 W=720e-9 AD=100.8e-15 AS=100.8e-15 PD=1.72e-6 PS=1.72e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i0__pm7 n6__r2 n8__i14__shift n8__i14__net2 n254__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i1__pm0 n9__i14__i1__net1 n9__i14__shift n258__vdd n254__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i1__pm5 n5__i14__net8 i14__i1__net1 n7__i14__net9 n254__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i1__pm7 n8__r1 n16__i14__shift n5__i14__net8 n254__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i2__pm0 n9__i14__i2__net1 n17__i14__shift n253__vdd n254__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i2__pm5 n4__i14__net14 i14__i2__net1 n7__i14__net15 n254__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i2__pm7 n11__r0 n24__i14__shift n4__i14__net14 n254__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i4__pm5 i14__i4__net1 n17__clkb i14__net15 n229__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i4__pm4 n252__vdd i14__i4__net5 i14__i4__net1 n229__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i4__pm2 i14__i4__net4 n2__i14__net8 n252__vdd n229__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i4__pm3 n6__i14__i4__net5 n21__clk i14__i4__net4 n229__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i5__pm1 n266__vdd n60__rst n5__i14__i5__rstb n229__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i5__pm0 n4__i14__i5__net5 i14__i5__rstb n266__vdd n229__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i5__pm5 i14__i5__net1 n21__clkb n6__serial_out n229__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i5__pm4 n268__vdd i14__i5__net5 i14__i5__net1 n229__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i5__pm2 i14__i5__net4 n2__i14__net14 n268__vdd n229__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i5__pm3 n6__i14__i5__net5 n25__clk i14__i5__net4 n229__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i3__pm4 n233__vdd i14__i3__net5 i14__i3__net1 n229__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i3__pm2 i14__i3__net4 n2__i14__net2 n233__vdd n229__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i3__pm3 n6__i14__i3__net5 n17__clk i14__i3__net4 n229__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i0__pm0 n9__i14__i0__net1 i14__shift n259__vdd n254__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i4__pm1 n249__vdd n54__rst n5__i14__i4__rstb n229__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i4__pm0 n4__i14__i4__net5 i14__i4__rstb n249__vdd n229__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i0__pm5 n8__i14__net2 i14__i0__net1 n219__vss n254__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i7__pm0 i14__i7__net2 n69__clk4 n264__vdd n261__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i7__pm1 n7__i14__i7__net1 n17__clk2 i14__i7__net2 n261__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i3__pm1 n228__vdd n48__rst n5__i14__i3__rstb n229__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i3__pm0 n4__i14__i3__net5 i14__i3__rstb n228__vdd n229__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i7__nm1 n28__i14__shift i14__i7__net1 n263__vdd n261__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i3__pm5 i14__i3__net1 n13__clkb i14__net9 n229__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi8__pm2 n2__i8__net49 n5__a2 n164__vdd n165__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi8__pm0 i8__net52 n7__a2 n159__vdd n165__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi8__pm3 n163__vdd a3 n2__i8__net49 n165__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi8__pm1 n8__i8__net51 n3__a3 i8__net52 n165__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi8__pm4 n9__s1 i8__net51 i8__net49 n165__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi8__pm5 n162__vdd i8__carry_bar n17__c1 n165__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi8__pm6 n4__i8__carry_bar n10__a2 n161__vdd n165__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi8__pm7 n152__vdd n6__a3 n4__i8__carry_bar n165__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi9__pm2 n2__i9__net49 s0 n203__vdd n180__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi9__pm0 i9__net52 n3__s0 n198__vdd n180__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi9__pm3 n202__vdd s1 n2__i9__net49 n180__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi9__pm1 n8__i9__net51 n3__s1 i9__net52 n180__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi9__pm4 r0 i9__net51 i9__net49 n180__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi9__pm5 n201__vdd i9__carry_bar n13__net12 n180__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi9__pm6 n4__i9__carry_bar n6__s0 n200__vdd n180__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi9__pm7 n191__vdd n6__s1 n4__i9__carry_bar n180__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi7__pm2 n2__i7__net49 n5__a0 n179__vdd n180__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi7__pm0 i7__net52 n7__a0 n174__vdd n180__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi7__pm3 n178__vdd a1 n2__i7__net49 n180__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi7__pm1 n8__i7__net51 n3__a1 i7__net52 n180__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi7__pm4 n9__s0 i7__net51 i7__net49 n180__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi7__pm5 n177__vdd i7__carry_bar n17__c0 n180__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi7__pm6 n4__i7__carry_bar n10__a0 n176__vdd n180__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi7__pm7 n167__vdd n6__a1 n4__i7__carry_bar n180__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi10__pm7 n220__vdd n9__c0 n7__i10__net122 n165__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi10__pm9 i10__net119 n9__net12 n11__i10__net114 n165__vdd g45p1svt L=45e-9 W=720e-9 AD=115.2e-15 AS=115.2e-15 PD=1.74e-6 PS=1.74e-6 NRD=1.16667 NRS=1.16667 M=1
mi10__pm10 i10__net118 n13__c1 i10__net119 n165__vdd g45p1svt L=45e-9 W=720e-9 AD=115.2e-15 AS=115.2e-15 PD=1.76e-6 PS=1.76e-6 NRD=1.16667 NRS=1.16667 M=1
mi10__pm11 n219__vdd n13__c0 i10__net118 n165__vdd g45p1svt L=45e-9 W=720e-9 AD=100.8e-15 AS=100.8e-15 PD=1.74e-6 PS=1.74e-6 NRD=1.16667 NRS=1.16667 M=1
mi10__pm12 r1 n2__i10__net114 n218__vdd n165__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi10__pm13 n4__r2 n5__i10__net116 n217__vdd n165__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi10__pm1 i10__net117 c0 n223__vdd n165__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi10__pm0 n13__i10__net116 c1 i10__net117 n165__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi10__pm2 n3__i10__net115 net12 n11__i10__net116 n165__vdd g45p1svt L=45e-9 W=960e-9 AD=153.6e-15 AS=153.6e-15 PD=2.22e-6 PS=2.22e-6 NRD=1.16667 NRS=1.16667 M=1
mi10__pm4 n222__vdd n5__c0 n3__i10__net115 n165__vdd g45p1svt L=45e-9 W=960e-9 AD=153.6e-15 AS=153.6e-15 PD=2.24e-6 PS=2.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi10__pm3 n7__i10__net115 n5__c1 n222__vdd n165__vdd g45p1svt L=45e-9 W=960e-9 AD=134.4e-15 AS=134.4e-15 PD=2.22e-6 PS=2.22e-6 NRD=1.16667 NRS=1.16667 M=1
mi10__pm5 n2__i10__net122 i10__net116 n7__i10__net114 n165__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi10__pm6 n221__vdd n5__net12 n2__i10__net122 n165__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi10__pm8 n7__i10__net122 n9__c1 n221__vdd n165__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi2__pm36 i2__net40 n22__clk4 n4__i2__net4 n109__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__pm35 n106__vdd n1__yin2 i2__net40 n109__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__pm33 i2__net12 i2__net4 n106__vdd n109__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__pm34 n17__y2 n21__clk4b i2__net12 n109__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__pm18 n4__i2__net2 n5__i2__rstb n105__vdd n109__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__pm26 i2__net28 n30__clk4 n4__i2__net2 n109__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__pm25 n104__vdd n1__yin3 i2__net28 n109__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__pm27 i2__net38 n2__i2__net2 n104__vdd n109__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__pm28 n19__y3 n33__clk4b i2__net38 n109__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__pm20 n96__vdd n8__i2__rstb n13__i2__net4 n109__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__pm16 n13__i2__rstb n21__rst n96__vdd n109__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__pm22 i2__net33 n6__clk4 n4__i2__net1 n109__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__pm21 n110__vdd n1__yin0 i2__net33 n109__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__pm24 i2__net35 n2__i2__net1 n110__vdd n109__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__pm23 n11__y0 n5__clk4b i2__net35 n109__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__pm17 n108__vdd i2__rstb n9__i2__net1 n109__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__pm19 n4__i2__net3 n3__i2__rstb n108__vdd n109__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__pm30 i2__net24 n14__clk4 n4__i2__net3 n109__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__pm29 n107__vdd n1__yin1 i2__net24 n109__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__pm31 i2__net26 n2__i2__net3 n107__vdd n109__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__pm32 n15__y1 n13__clk4b i2__net26 n109__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__pm36 i1__net40 n24__clk4 n4__i1__net4 n124__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__pm35 n121__vdd n1__xin2 i1__net40 n124__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__pm33 i1__net12 i1__net4 n121__vdd n124__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__pm34 n17__x2 n23__clk4b i1__net12 n124__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__pm18 n4__i1__net2 n5__i1__rstb n120__vdd n124__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__pm26 i1__net28 n32__clk4 n4__i1__net2 n124__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__pm25 n119__vdd n1__xin3 i1__net28 n124__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__pm27 i1__net38 n2__i1__net2 n119__vdd n124__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__pm28 n19__x3 n35__clk4b i1__net38 n124__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__pm20 n111__vdd n8__i1__rstb n13__i1__net4 n124__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__pm16 n13__i1__rstb n25__rst n111__vdd n124__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__pm22 i1__net33 n8__clk4 n4__i1__net1 n124__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__pm21 n125__vdd n1__xin0 i1__net33 n124__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__pm24 i1__net35 n2__i1__net1 n125__vdd n124__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__pm23 n14__x0 n7__clk4b i1__net35 n124__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__pm17 n123__vdd i1__rstb n9__i1__net1 n124__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__pm19 n4__i1__net3 n3__i1__rstb n123__vdd n124__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__pm30 i1__net24 n16__clk4 n4__i1__net3 n124__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__pm29 n122__vdd n1__xin1 i1__net24 n124__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__pm31 i1__net26 n2__i1__net3 n122__vdd n124__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__pm32 n15__x1 n15__clk4b i1__net26 n124__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__pm30 n133__vdd i0__net4 i0__net20 n124__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__pm31 i0__net13 n2__i0__net6 n133__vdd n124__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__pm32 n7__i0__net3 n6__i0__net1 i0__net13 n124__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__pm33 n14__i0__net4 i0__net3 n130__vdd n124__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__pm34 n33__clk4 n4__i0__net4 n128__vdd n124__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__pm35 n29__clk4b clk4 n131__vdd n124__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__pm23 i0__net16 n2__clk n4__i0__net2 n124__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__pm22 n137__vdd i0__net1 i0__net16 n124__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__pm24 i0__net19 n2__i0__net2 n137__vdd n124__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__pm25 n11__clk2 n3__clkb i0__net19 n124__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__pm26 n14__i0__net1 clk2 n136__vdd n124__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__pm29 i0__net20 n6__clk2 n4__i0__net6 n124__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi11__pm0 n274__vdd n3__serial_out n3__i11__net1 n272__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi12__m4_99__rcx n390__vss n344__i12__net3 n383__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_98__rcx n391__r_out n347__i12__net3 n390__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_97__rcx n392__vss n350__i12__net3 n391__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_96__rcx n399__r_out n353__i12__net3 n392__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_95__rcx n394__vss n356__i12__net3 n399__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_94__rcx n403__r_out n359__i12__net3 n394__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=699.75e-15 AS=699.75e-15 PD=9.68e-6 PS=9.68e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_93__rcx n384__vss n326__i12__net3 n359__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_92__rcx n367__r_out n329__i12__net3 n384__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_91__rcx n386__vss n332__i12__net3 n367__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_90__rcx n375__r_out n335__i12__net3 n386__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_89__rcx n388__vss n338__i12__net3 n375__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_88__rcx n383__r_out n341__i12__net3 n388__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_87__rcx n359__r_out n323__i12__net3 n382__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_86__rcx n335__r_out n305__i12__net3 n376__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_85__rcx n378__vss n308__i12__net3 n335__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_84__rcx n343__r_out n311__i12__net3 n378__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_83__rcx n380__vss n314__i12__net3 n343__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_82__rcx n351__r_out n317__i12__net3 n380__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_81__rcx n382__vss n320__i12__net3 n351__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_80__rcx n311__r_out n287__i12__net3 n370__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_79__rcx n372__vss n290__i12__net3 n311__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_78__rcx n319__r_out n293__i12__net3 n372__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_77__rcx n374__vss n296__i12__net3 n319__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_76__rcx n327__r_out n299__i12__net3 n374__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_75__rcx n376__vss n302__i12__net3 n327__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_74__rcx n287__r_out n269__i12__net3 n364__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_73__rcx n366__vss n272__i12__net3 n287__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_72__rcx n295__r_out n275__i12__net3 n366__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_71__rcx n368__vss n278__i12__net3 n295__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_70__rcx n303__r_out n281__i12__net3 n368__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_69__rcx n370__vss n284__i12__net3 n303__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_68__rcx n263__r_out n251__i12__net3 n358__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_67__rcx n360__vss n254__i12__net3 n263__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_66__rcx n271__r_out n257__i12__net3 n360__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_65__rcx n362__vss n260__i12__net3 n271__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_64__rcx n279__r_out n263__i12__net3 n362__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_63__rcx n364__vss n266__i12__net3 n279__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_62__rcx n358__vss n248__i12__net3 n255__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_61__rcx n352__vss n230__i12__net3 n231__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_60__rcx n239__r_out n233__i12__net3 n352__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_59__rcx n354__vss n236__i12__net3 n239__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_58__rcx n247__r_out n239__i12__net3 n354__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_57__rcx n356__vss n242__i12__net3 n247__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_56__rcx n255__r_out n245__i12__net3 n356__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_55__rcx n346__vss n212__i12__net3 n207__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_54__rcx n215__r_out n215__i12__net3 n346__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_53__rcx n348__vss n218__i12__net3 n215__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_52__rcx n223__r_out n221__i12__net3 n348__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_51__rcx n350__vss n224__i12__net3 n223__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_50__rcx n231__r_out n227__i12__net3 n350__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_49__rcx n340__vss n194__i12__net3 n179__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_48__rcx n191__r_out n197__i12__net3 n340__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_47__rcx n342__vss n200__i12__net3 n191__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_46__rcx n199__r_out n203__i12__net3 n342__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_45__rcx n344__vss n206__i12__net3 n199__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_44__rcx n207__r_out n209__i12__net3 n344__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_43__rcx n333__vss n176__i12__net3 n159__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_42__rcx n167__r_out n179__i12__net3 n333__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_41__rcx n335__vss n182__i12__net3 n167__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_40__rcx n175__r_out n185__i12__net3 n335__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_39__rcx n337__vss n188__i12__net3 n175__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_38__rcx n179__r_out n191__i12__net3 n337__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_37__rcx n159__r_out n173__i12__net3 n331__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_36__rcx n135__r_out n155__i12__net3 n325__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_35__rcx n327__vss n158__i12__net3 n135__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_34__rcx n143__r_out n161__i12__net3 n327__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_33__rcx n329__vss n164__i12__net3 n143__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_32__rcx n151__r_out n167__i12__net3 n329__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_31__rcx n331__vss n170__i12__net3 n151__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_30__rcx n111__r_out n137__i12__net3 n319__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_29__rcx n321__vss n140__i12__net3 n111__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_28__rcx n119__r_out n143__i12__net3 n321__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_27__rcx n323__vss n146__i12__net3 n119__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_26__rcx n127__r_out n149__i12__net3 n323__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_25__rcx n325__vss n152__i12__net3 n127__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_24__rcx n87__r_out n119__i12__net3 n313__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_23__rcx n315__vss n122__i12__net3 n87__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_22__rcx n95__r_out n125__i12__net3 n315__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_21__rcx n317__vss n128__i12__net3 n95__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_20__rcx n103__r_out n131__i12__net3 n317__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_19__rcx n319__vss n134__i12__net3 n103__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_18__rcx n63__r_out n101__i12__net3 n307__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_17__rcx n309__vss n104__i12__net3 n63__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_16__rcx n71__r_out n107__i12__net3 n309__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_15__rcx n311__vss n110__i12__net3 n71__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_14__rcx n79__r_out n113__i12__net3 n311__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_13__rcx n313__vss n116__i12__net3 n79__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_12__rcx n307__vss n88__i12__net3 n55__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_11__rcx n301__vss n40__i12__net3 n31__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_10__rcx n39__r_out n53__i12__net3 n301__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_9__rcx n303__vss n56__i12__net3 n39__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_8__rcx n47__r_out n69__i12__net3 n303__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_7__rcx n305__vss n72__i12__net3 n47__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_6__rcx n55__r_out n85__i12__net3 n305__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_5__rcx n15__r_out n5__i12__net3 n295__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_4__rcx n297__vss n8__i12__net3 n15__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_3__rcx n23__r_out n21__i12__net3 n297__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_2__rcx n299__vss n24__i12__net3 n23__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4_1__rcx n31__r_out n37__i12__net3 n299__vss n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.73e-6 PS=9.73e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m4 n295__vss n2__i12__net3 n7__r_out n7__vss g45n2svt L=150e-9 W=4.665e-6 AD=933e-15 AS=933e-15 PD=9.68e-6 PS=9.68e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m3_10__rcx n50__i12__net3 n14__i12__net2 n276__vss n7__vss g45n2svt L=150e-9 W=4.715e-6 AD=943e-15 AS=943e-15 PD=9.83e-6 PS=9.83e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m3_9__rcx n280__vss n17__i12__net2 n50__i12__net3 n7__vss g45n2svt L=150e-9 W=4.715e-6 AD=943e-15 AS=943e-15 PD=9.83e-6 PS=9.83e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m3_8__rcx n66__i12__net3 n20__i12__net2 n280__vss n7__vss g45n2svt L=150e-9 W=4.715e-6 AD=943e-15 AS=943e-15 PD=9.83e-6 PS=9.83e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m3_7__rcx n284__vss n23__i12__net2 n66__i12__net3 n7__vss g45n2svt L=150e-9 W=4.715e-6 AD=943e-15 AS=943e-15 PD=9.83e-6 PS=9.83e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m3_6__rcx n82__i12__net3 n26__i12__net2 n284__vss n7__vss g45n2svt L=150e-9 W=4.715e-6 AD=943e-15 AS=943e-15 PD=9.83e-6 PS=9.83e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m3_5__rcx n288__vss n29__i12__net2 n82__i12__net3 n7__vss g45n2svt L=150e-9 W=4.715e-6 AD=943e-15 AS=943e-15 PD=9.83e-6 PS=9.83e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m3_4__rcx n366__i12__net3 n39__i12__net2 n288__vss n7__vss g45n2svt L=150e-9 W=4.715e-6 AD=707.25e-15 AS=707.25e-15 PD=9.78e-6 PS=9.78e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi11__m0 n254__vss n2__serial_out n4__net5 n7__vss g45n2svt L=150e-9 W=2.32e-6 AD=464e-15 AS=464e-15 PD=4.99e-6 PS=4.99e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi11__m3 n9__r_in n2__i11__net1 n254__vss n7__vss g45n2svt L=150e-9 W=2.32e-6 AD=348e-15 AS=348e-15 PD=4.99e-6 PS=4.99e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m7 n9__i12__net1 n4__r_in n267__vss n7__vss g45n2svt L=150e-9 W=640e-9 AD=96e-15 AS=96e-15 PD=1.58e-6 PS=1.58e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m0_1__rcx n269__vss n2__i12__net1 n36__i12__net2 n7__vss g45n2svt L=150e-9 W=2.88e-6 AD=576e-15 AS=576e-15 PD=6.11e-6 PS=6.11e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m0 n47__i12__net2 n5__i12__net1 n269__vss n7__vss g45n2svt L=150e-9 W=2.88e-6 AD=432e-15 AS=432e-15 PD=6.11e-6 PS=6.11e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m3_3__rcx n18__i12__net3 n2__i12__net2 n258__vss n7__vss g45n2svt L=150e-9 W=4.715e-6 AD=943e-15 AS=943e-15 PD=9.78e-6 PS=9.78e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m3_2__rcx n272__vss n5__i12__net2 n18__i12__net3 n7__vss g45n2svt L=150e-9 W=4.715e-6 AD=943e-15 AS=943e-15 PD=9.83e-6 PS=9.83e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m3_1__rcx n34__i12__net3 n8__i12__net2 n272__vss n7__vss g45n2svt L=150e-9 W=4.715e-6 AD=943e-15 AS=943e-15 PD=9.83e-6 PS=9.83e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi12__m3 n276__vss n11__i12__net2 n34__i12__net3 n7__vss g45n2svt L=150e-9 W=4.715e-6 AD=943e-15 AS=943e-15 PD=9.83e-6 PS=9.83e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi6__nm0 n72__vss n3__x3 n6__i6__abar n7__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi6__nm1 n6__i6__bbar n3__y3 n72__vss n7__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi6__nm2 n11__a3 n7__x3 n2__i6__net3 n7__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi6__nm4 i6__net4 n3__i6__bbar n11__a3 n7__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi6__nm5 n77__vss n3__i6__abar i6__net4 n7__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi6__nm3 i6__net3 n7__y3 n77__vss n7__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__nm0 n73__vss n3__x2 n6__i5__abar n7__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__nm1 n6__i5__bbar n3__y2 n73__vss n7__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__nm2 n3__a2 n7__x2 n2__i5__net3 n7__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__nm4 i5__net4 n3__i5__bbar n3__a2 n7__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__nm5 n44__vss n3__i5__abar i5__net4 n7__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__nm3 i5__net3 n7__y2 n44__vss n7__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi4__nm0 n76__vss n3__x1 n6__i4__abar n7__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi4__nm1 n6__i4__bbar n3__y1 n76__vss n7__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi4__nm2 n11__a1 n7__x1 n2__i4__net3 n7__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi4__nm4 i4__net4 n3__i4__bbar n11__a1 n7__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi4__nm5 n118__vss n3__i4__abar i4__net4 n7__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi4__nm3 i4__net3 n10__y1 n118__vss n7__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi3__nm0 n43__vss n3__x0 n6__i3__abar n7__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi3__nm1 n6__i3__bbar n3__y0 n43__vss n7__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi3__nm2 n3__a0 n7__x0 n2__i3__net3 n7__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi3__nm4 i3__net4 n3__i3__bbar n3__a0 n7__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi3__nm5 n46__vss n3__i3__abar i3__net4 n7__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi3__nm3 i3__net3 n7__y0 n46__vss n7__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi15__nm0 n8__clkb n6__clk n5__vss n7__vss g45n1svt L=45e-9 W=360e-9 AD=50.4e-15 AS=50.4e-15 PD=1e-6 PS=1e-6 NRD=1.16667 NRS=1.16667 M=1
mi14__i0__nm8 n8__r2 n3__i14__i0__net1 n9__i14__net2 n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i1__nm0 n6__i14__i1__net1 n12__i14__shift n248__vss n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i1__nm6 n7__i14__net8 n13__i14__shift n9__i14__net9 n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i1__nm8 n10__r1 n3__i14__i1__net1 n7__i14__net8 n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i2__nm0 n7__i14__i2__net1 n20__i14__shift n249__vss n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i2__nm6 n6__i14__net14 n21__i14__shift n9__i14__net15 n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i2__nm8 n10__r0 n3__i14__i2__net1 n6__i14__net14 n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i4__nm3 i14__i4__net2 n20__clk n3__i14__net15 n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i4__nm4 n234__vss n3__i14__i4__net5 i14__i4__net2 n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i4__nm2 i14__i4__net3 n3__i14__net8 n234__vss n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i4__nm1 n8__i14__i4__net5 n18__clkb i14__i4__net3 n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i5__nm0 n233__vss n59__rst n4__i14__i5__rstb n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i5__nm16 n10__serial_out n62__rst n233__vss n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i5__nm3 i14__i5__net2 n24__clk n8__serial_out n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i5__nm4 n223__vss n3__i14__i5__net5 i14__i5__net2 n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i5__nm2 i14__i5__net3 n3__i14__net14 n223__vss n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i5__nm1 n8__i14__i5__net5 n22__clkb i14__i5__net3 n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i3__nm4 n236__vss n3__i14__i3__net5 i14__i3__net2 n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i3__nm2 i14__i3__net3 n3__i14__net2 n236__vss n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i3__nm1 n8__i14__i3__net5 n14__clkb i14__i3__net3 n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i0__nm0 n7__i14__i0__net1 n4__i14__shift n246__vss n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i4__nm0 n235__vss n53__rst n4__i14__i4__rstb n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i4__nm16 n5__i14__net15 n56__rst n235__vss n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i0__nm6 n9__i14__net2 n5__i14__shift n217__vss n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i7__nm4 n5__i14__i7__net1 n71__clk4 n240__vss n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i7__nm5 n242__vss n19__clk2 n5__i14__i7__net1 n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i3__nm0 n237__vss n47__rst n4__i14__i3__rstb n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i3__nm16 n5__i14__net9 n50__rst n237__vss n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i7__nm0 n27__i14__shift n4__i14__i7__net1 n244__vss n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi14__i3__nm3 i14__i3__net2 n16__clk n3__i14__net9 n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi8__nm3 i8__net50 n8__a2 n12__s1 n7__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi8__nm0 n5__i8__net51 n9__a2 n150__vss n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi8__nm4 n149__vss n4__a3 i8__net50 n7__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi8__nm1 n147__vss n5__a3 n5__i8__net51 n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi8__nm2 n146__vss n3__i8__net51 n13__s1 n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi8__nm5 n145__vss n3__i8__carry_bar n19__c1 n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi8__nm7 i8__net1 n12__a2 n6__i8__carry_bar n7__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi8__nm6 n139__vss n8__a3 i8__net1 n7__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi9__nm3 i9__net50 n4__s0 n4__r0 n7__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi9__nm0 n5__i9__net51 n5__s0 n186__vss n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi9__nm4 n185__vss n4__s1 i9__net50 n7__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi9__nm1 n183__vss n5__s1 n5__i9__net51 n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi9__nm2 n182__vss n3__i9__net51 n5__r0 n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi9__nm5 n181__vss n3__i9__carry_bar n16__net12 n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi9__nm7 i9__net1 n8__s0 n6__i9__carry_bar n7__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi9__nm6 n169__vss n8__s1 i9__net1 n7__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi7__nm3 i7__net50 n8__a0 n12__s0 n7__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi7__nm0 n5__i7__net51 n9__a0 n193__vss n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi7__nm4 n192__vss n4__a1 i7__net50 n7__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi7__nm1 n190__vss n5__a1 n5__i7__net51 n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi7__nm2 n189__vss n3__i7__net51 n13__s0 n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi7__nm5 n188__vss n3__i7__carry_bar n20__c0 n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi7__nm7 i7__net1 n12__a0 n6__i7__carry_bar n7__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi7__nm6 n187__vss n8__a1 i7__net1 n7__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi10__nm6 n205__vss n12__c0 n5__i10__net125 n7__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi10__nm11 i10__net120 n12__net12 n13__i10__net114 n7__vss g45n1svt L=45e-9 W=360e-9 AD=57.6e-15 AS=57.6e-15 PD=1.02e-6 PS=1.02e-6 NRD=1.16667 NRS=1.16667 M=1
mi10__nm9 i10__net121 n16__c1 i10__net120 n7__vss g45n1svt L=45e-9 W=360e-9 AD=57.6e-15 AS=57.6e-15 PD=1.04e-6 PS=1.04e-6 NRD=1.16667 NRS=1.16667 M=1
mi10__nm10 n204__vss n16__c0 i10__net121 n7__vss g45n1svt L=45e-9 W=360e-9 AD=50.4e-15 AS=50.4e-15 PD=1.02e-6 PS=1.02e-6 NRD=1.16667 NRS=1.16667 M=1
mi10__nm12 n3__r1 n3__i10__net114 n203__vss n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi10__nm13 n3__r2 n8__i10__net116 n194__vss n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi10__nm0 i10__net123 n4__c0 n208__vss n7__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi10__nm1 n17__i10__net116 n4__c1 i10__net123 n7__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi10__nm2 n3__i10__net124 n4__net12 n14__i10__net116 n7__vss g45n1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi10__nm3 n207__vss n8__c0 n3__i10__net124 n7__vss g45n1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi10__nm4 n8__i10__net124 n8__c1 n207__vss n7__vss g45n1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi10__nm8 n2__i10__net125 n4__i10__net116 n10__i10__net114 n7__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi10__nm5 n206__vss n8__net12 n2__i10__net125 n7__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi10__nm7 n5__i10__net125 n12__c1 n206__vss n7__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm38 i2__net41 n18__clk4b n7__i2__net4 n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm39 n89__vss n3__yin2 i2__net41 n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm37 i2__net13 n2__i2__net4 n89__vss n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm36 n15__y2 n25__clk4 i2__net13 n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm18 n88__vss n9__rst n15__y2 n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm46 i2__net37 n26__clk4b n7__i2__net2 n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm47 n87__vss n3__yin3 i2__net37 n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm45 i2__net39 n3__i2__net2 n87__vss n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm44 n17__y3 n37__clk4 i2__net39 n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm17 n79__vss n13__rst n16__y3 n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm35 n16__i2__rstb n24__rst n79__vss n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm48 i2__net34 n2__clk4b n7__i2__net1 n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm49 n92__vss n3__yin0 i2__net34 n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm51 i2__net36 n3__i2__net1 n92__vss n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm50 n13__y0 n9__clk4 i2__net36 n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm16 n91__vss n1__rst n13__y0 n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm19 n4__y1 n6__rst n91__vss n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm42 i2__net25 n10__clk4b n7__i2__net3 n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm43 n90__vss n3__yin1 i2__net25 n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm41 i2__net27 n3__i2__net3 n90__vss n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm40 n16__y1 n17__clk4 i2__net27 n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm38 i1__net41 n20__clk4b n7__i1__net4 n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm39 n109__vss n3__xin2 i1__net41 n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm37 i1__net13 n2__i1__net4 n109__vss n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm36 n15__x2 n27__clk4 i1__net13 n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm18 n108__vss n11__rst n15__x2 n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm46 i1__net37 n28__clk4b n7__i1__net2 n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm47 n107__vss n3__xin3 i1__net37 n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm45 i1__net39 n3__i1__net2 n107__vss n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm44 n17__x3 n39__clk4 i1__net39 n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm17 n93__vss n15__rst n16__x3 n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm35 n16__i1__rstb n28__rst n93__vss n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm48 i1__net34 n4__clk4b n7__i1__net1 n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm49 n112__vss n3__xin0 i1__net34 n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm51 i1__net36 n3__i1__net1 n112__vss n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm50 n16__x0 n11__clk4 i1__net36 n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm16 n111__vss n3__rst n16__x0 n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm19 n8__x1 n8__rst n111__vss n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm42 i1__net25 n12__clk4b n7__i1__net3 n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm43 n110__vss n3__xin1 i1__net25 n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm41 i1__net27 n3__i1__net3 n110__vss n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__nm40 n16__x1 n19__clk4 i1__net27 n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__nm17 n116__vss n3__i0__net4 i0__net34 n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__nm18 i0__net15 n3__i0__net6 n116__vss n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__nm19 n6__i0__net3 n7__clk2 i0__net15 n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__nm21 n12__i0__net4 n4__i0__net3 n115__vss n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__nm23 n36__clk4 n7__i0__net4 n113__vss n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__nm22 n30__clk4b n4__clk4 n114__vss n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__nm10 i0__net17 n2__clkb n7__i0__net2 n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__nm11 n106__vss n3__i0__net1 i0__net17 n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__nm12 i0__net33 n3__i0__net2 n106__vss n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__nm13 n12__clk2 n7__clk i0__net33 n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__nm14 n12__i0__net1 n4__clk2 n117__vss n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi0__nm20 i0__net34 n5__i0__net1 n7__i0__net6 n7__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi11__nm0 n252__vss n5__serial_out n6__i11__net1 n7__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
.ENDS PIPO_and_Combinational
